// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
kXjW0mtn1GvZH8QKJ4WfklrA8qKWG0lu4ZWHct3yWJXraV+JnFz6y9aigDn18ut2MBdteC4NRiNP
CrnStIJsfprr8SwH9MzWB+l2bIEwUpkuK3yTPVCoXUhlZrIi58W+3QyLNVTBzqUA3uSwP68FdAWt
h1xBu+4LL4QCUQU/bQvDskj+mrBwdVgmrTYeaJ5Zjzvjyk9RVPMZDdduSH+ou614aJ5CfJr47/XH
Lv0DLB6HzJ3XWz67AAAj0pEg08cxz7lGPxsQ9G4UWvtR5z5ZsAVydFFnZ2KnAaNDymC4HLU/uvEH
A3CQ+vpfnYmdVdsMqfPZd2qLy/UhEM+wtG0ACA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5104)
AXovTvj4piXWhyfgfqKW3+8MkQdioi+OelFcNTsI0Q5D8CqbAkZNt396s9+A8HDgiUJuZD8kH7iR
ao8vbYUGc+XjxY/WkOQlNLFDcFVKeX9Q2r0NxQkdtna3tGxThezhiT7iti9zhGkpw9nKezgJFVpE
bwqLAUWsKKlPNJpvEVpDExWV2HvPMEPFgrQ4Ln9jYKIyybiRWm2jFiwMAcHwB2mv5XjereyutWQO
EwrF9MzYBQ0St270GX+uO0UQAUk+9TMHant7WvESazsGHLRpnigV45G/8epHjuiDtHXF+lZ81E8B
sJjofPizYKaEifD3MKS/PaXVIIsIENkwBvWIFWMurbrik0Hjgc0UaJLc1XO5UDTV71AG6yp6nNPf
Cd10jmo/Ybyv3WkY8+fBeoV51X9JwN0+Pb3H6vHV3j5XwTd+4baqg2TvQvHucebQ7XvsAj6fCNXv
XhVr1SfYNGcgsus/9fUkWCNEn7ak/qQtv9a/cvyfnOsG9ZipXhl5Gg+AE09mB7A8U3VITbOia9+q
adOI3D3KtvVTPyavLOQk8JgYlqPaK05tJhcuC2AqR/WhrPgkX8h6hfeVo7HK4cEcATJ1Kqf7l8Yn
asLvmiGO5oGPFBLOs6bw+UM5EO9iU0+ld0NDptGZshIwDM3o0Y5Uv7B9SZqH9e/toWGAU/jVE/mQ
+z0tyx/i9LqqyiokghHJ7S0qhuxlYyJNUMEoRhAXSNLYcQYcqRh985Y5TDUE1eCNHuGQx5Q0oXKJ
e6+9zDZFWVe2O30+s6uPLFZnM1BlZVwyUCKHGItpGKVEXJvQTbRvIQ11iLV2A9VFhtLB3JhWAnQi
Qrtl2j6phgvQQwP9fdoO3nciwRe26QZCJ4WBfmxy8QYG548fAAhU3rV07cetxRkRRYETZJEBn8Kd
p1s2UkZqOXrwMAZKwjpGTeS/PX8rUJcuYPMiMnc0w1zd6alptUz1RCHkI0mbHnuAgn2ev84EYGyl
/SzEsL7o7Y6cBEb27tjM07afscFlAmN86N/jc8m+ufAqE1JfU5iFrFJyILiZt+hTSn75Tfn6rmZ0
Tn08caodMdYf2p9fM4HOoNGJFYwm41aufVeVQeAGO6tYiMYiI6t3KlfyXDoDYpzQeb3fWljzale3
tA06gJ9kMK8Rkmkfk4SRsV3CfSbeMGEh0rxMVpzFs81dtNigmatSg/ObQtj4+VPg/6E5QXOAI7bC
hpOyho9GotZhMgq+nrGqErBD2gtOyNJUHyzkZijxCxR7vFuPi3pDyDThvhMO4rOjGISQ+o1fKllx
ef46fbUrlZAsjJ1wRKbnnymD9go6Giy8IIiMCXIYsBA2gh38WFfLW+szgT4Fk3DA8301Rw1Gh4oy
Uf25R3AhSmds6Mwr1JMHdNtRrWIiN08UZ3122BAZyl7ccpH/AlLb06KZtUl0WRqaZ4ma7EfgRhk+
pRkWafkmhVJANgBBq89ZgCK7/qBsSyNR9mpKXAPQNDlzmgvT0ng8PcNUBUCFP1fdm1e0ENb0bUOf
V97G0rvrX6DquY+l8vdx8rW0EZ6HxgWniIjy7WsVqc/z5wxoMTdNES0a+RWkknwseBUIFVRo9I6g
DTwdhPIATnokzEAO4KthAmpdHkU9En3vRNHJvy6pvU9WUo1Ny8x3dnvPgdF00+atZDYrtXnPmEUz
YzDeOOikT9RJCJ2OIbclNW6V6amVd3/OQgcetvzY63KLnt/+kj/xcmWBYUrutQx5iLeAggY3WZxq
YdDdFYvI5voyUWZBTTuQ3ifIDexP5BZFlgL9gRu2TzNc0bwZpmMFHs5kKChze5pgP6N5LF72QKBp
zM54gLNt66nSqPfTSr41aGr9DMthKHvv0nhiXSCy2h9ed0c7vfyjcfz7dg7kbVQxOsk7trnpdIiq
kjF6cIq5mPDtcU5bHt+TEMb1MlkDnVgHGf8GOVn9FBS3GcS+ThQ2KPxHjq/ebaNm3peeqNQAeodw
F9UIdKEU4OUxkFoWsELQuYK9V8rPSuxZZEpQ3U04EGJiBvYJcp2wCfCs5NwahOz8TBU/xhTbNshb
5mm+S1cJAB08JSEkrVUL5lVu0+EQEazWOh+CwYkWxCdCY0RbeVISZ2HZTUBLZ3Dd3N9TzX7o+Tat
HNsfHFB106s8xjPwYlAJD8Tk4r0vCaQyaMYagdqzPI5e65d+/AaHIcfT7JD2hSGOMiydYEqNI0/l
ww+zk71w6l0AgiFoWIvIK1h5Tpb4GQKgwLHEgXqhfyYQAQj0EEJ72d95yLvAX/E2Vmfbh771f7tF
U9Gm+Llmi4Nz/YjuGAoNVUJSqGrcYAUUQTNpbjtGnTsCgZWWlm/AYfxuXXJn9YXAcFXzKN3ZBRBH
iP1yuqoPcOsfM4WQEtebTqRSVC+elY7km+HoGUN0cDyTM6qo03EqS070BmfJqkl8g1rY6XEV5YVH
bj7kcCGVk89jPYRxnzk9ijpz18BV3d5el0SYf3vyqYMP7/wwYmDvid/QzSnOnSxfNn5s6Pm/Yshd
o97fyp5DY4kHaMKM2DHZQJbgta6UaOeZTnO6R3afHRbvuGNubdHzmLv2bXTGiwFI/QpkF+BJ/S3Y
WMLOp00wJFWxfsmLr3wvHDiZ+3RSXWIY7Xq524ZCvkce6JELZI7fgBGta4JGKJNl10KaMj9aZCbL
pxdgzsbiskTkvKISyhtdEz/OLDE5BQcKGk7XLqzRtMr4CF6ewoDUM0TRSW80avKVvYXPDftBwUwi
1IGbvHq4C6w7A7K/U3Og6lWHnOQlmlQgvB8u/BDvwVy254LpMB7lh1a50IlFY8jXJapTWIXNPyDP
vh4olXFjJVB20aTsjQJI3plsv74I/V3rO/OwSQbhm5IPaBhM79ENZpz80Y15icgCTVLKzmd9Pi9C
HZD0cgY4DWZigZaL84fc61EizkcF+dEXlu/KBFrDxH5QVkVtguOTZnbFhw+JKnqGG5veHXs+ZgpQ
OzF3RsgPazhXDyJknsiZWMXjcj0rWJgW2iNcRfD0Qd6YHtaDMfOEcs+7665c2+4ZUUZfAYslnbW8
4QT4KM8dNOGRLJeEDeyweCWFSM+b78VC0dYSDBEGMnyh9r8DnceU7eXAVgO3JkyecpOUk/STtYhV
WGj4Jrmr1aRZZ1AqKR6ShNa/ObPf26A1schUYurbmlDvbmKISv+LSux4juoB3QoPOr32bNvQNh4Y
KUEOR3i54REG1KHLwLcmZzmGV2e292TgXbtbP42QuFO3S00IqKt9aZBbhkESDbrW5/6TYYlTaNL8
J7OgTo3jpTpwt6ZKPXOl/HtHy0kh3KtAd+yvnYpDkb9PazHnmNZq8R7XQ61aEihOwoJxhLQ7SNs8
WcKM1u77nrHyzwFbST9jeonUYHq1WXMKWVW3/EWv7ebOVi3qkmaPUAx50WxD+7oPrPGFcOXq1QJ9
rowT2nLn3/iIWtMaXE5lVP6HKY38Oy1PrqJU2Uus3KY0bS6hE8eZDW3XU3xuVpFvcZtADghBhSLO
Q13oP4lDs0UqfM79NgWWgbZk49iM/F4DMd1PJvksSB53x6xofgtFHvYbWLsIlF6kt3WQK4ld7R0S
gzPjgx4uNeZ4mRJ1LxoysoLTZsQ0pdmQUwjqfWtzMyJpePtd1jeHvTgJC5T3euwdQQ5455Fs24r3
HBoYTwdWJVTtqx/spAkZo5adXwdLhnLZrDYkojD8yjD6aRgDKgz/CVZdKfzX3o0AWZ21ohV1WGRq
XyjUji2LNpinjKlse34hVrJZaxOc23N/MQ3Z0v7+kVBPJL9tymBoMoSEqhmkix4uOUwomgtUyw5H
YCgeDCcJUits0HTQ3Jtq/+NTiwxq2G3cFcF09hp9/8cu0x71I7jyrqXxglPAKvc2jTb0TmAry69P
QQp7DUMg3vwvG4lh6Z0ETFV0NUb/omEVX+7yRSEVx1ut6ozJ9dXv2jZyER2ea1KOmYsZrCpsG0MI
AQAAykv85eRutRIc6SYx0nU6A4MC/IQ/Md5lwNfQy6WGmtr7RxeP9ju3Ib8hBX+8o5mJ0sev/P4d
/ZEOUxNAz+jrVpZbn5t9tANERNWXPZVxWVtOOf5WEHRcF1gaQekb2jP2RyXUsXiPwQQiZgYF4HID
DDnAvYkWh+AQSZlwn62updmYtrB24Ln+zC014bRsPFDQvxd5Q9moGUQiKU+DB3SKO4rFtgmyAy+n
ARg1QXyuc7IpOEuKE2G6OS37XwzLLqa2ypW1Z1h7XUgmKT69dfEcUjuJ5yiOFGj7ho10+pkxjkuQ
8BurHjoebGfeHN7CziJVsxbggnQonIGCIrabEZOQbf7K0RkS+OoB0f4g/cDOwSjO/WwCyrKySQmB
EMNokVbXcFobZ8apc48Zr9i6kEGQEALiTZcP6xL545+lOpCILBE0MYWwdwJQmUFqwOJtbKs4huuM
WY/NhDwAMjCNjtGtevvFnCJl0yqpVmqnB1nm0FYjLoj6xM/3DimND75432aNdvMaRnbont/xxCt6
iQkxzz2+ovOfTk5oIrL6TUf0zy6dym3hWerBcA4GC48cLS19boFQA9PEcegK6PSO/rnI+LyUDidL
mikPP2my8wcEiekvM520qiNGP51wMXACP24d7/78AWTDCH6pQGM+1MSsv8s0ao3sr7gQ1mhsecSb
dZubYuZThhyWeDWCPLjdgEXTCZRx2+SoFk5q2hsgfOBbW40drab95IthUqZTgP58Bua0kOu5eR23
12nSO9fwEB0FgAnLhqm9+VuNkvABn/UKhs3tlyXKQIAaDhgRTpaSXpInKNk7FS/RZIQkV1afpKBh
z2gS3dnnCWMRTO4CHmREgYPngaA+s+I1l+4VOJbnwb5zYJN+RP1iQqc1jbR2GOgT6c2gEMxjt70W
HBEfxmafkx3cHjAMcEE9U4zBOKCT59vvLUCxi0Z11AopGLSXNSgkdSkQS2LjDmLD7/MslhgcAHGc
myhKyGdabLbmGyL4U2+nXFZkOoDmQsm2Q4UzeejR2Fg0p7L+airg672CXix1RwE8wXMJ0hRrBYVn
SqxTh8KpJohduwzzZLe462oE5yhvKIWuA0CG+7FnddHFkxB1dgt0cL2h3gnig84QZoQO8q2Zizso
+vfokrxFujBNg7jfFrSPHHf+eJsPcPr2UcTu3us2tf9akl0HKVoifKf3peOn8qEOXrGjDwutPVSK
k5ij00fSQdwdSo4pgGhtYPv21DCSHwLnq4XCk4PyQDAQQkOH7x9nZhAN2Y9EpxkMC/ZJ5bXjGLOs
kefPSThzhSHD3ddNk9IuUVhE2bjyru8pTjyuGYPEHBFq7aNML7QD8i1GFmIkWbQercd9WlWGOXOc
d7iN23Barj4bOkEOdrIatKLT2gYFHndApP/EFDpmc5rSWJS1c4GUc0s69GVNxT2QdptpWA4IJRCE
nDBseKCWx9Llq5St/K4fS8pzduYxso6jfWD2QZasQLW1uLXVXp4LDiXCosuT9EO4kd7wRpNfxmQl
Evz7l/U8VmrODXHXhZL61YsT9sjrlbIIXBe/qNSWT8RF4zGMuC7B0wLKZEoNMv/74zui3b6+n5XK
CdGM1YL3AKzCjgoI22tQSP/eHggMZamI2uh+l6jDjNbe2jXOhzCe/bLxEKfeIcZXZPo/CB6XScZy
1BB7QfwJDC7e7srKZOtiKqcY4iuf5OH1NRgB+H9qNnbxIu78MIY793xeIn97Ud3uKTt4BXOirMhI
0D8rvhnAfZgFYYNS/FlLfSUfP9tReswBPFF2JwxwpL/shCegt54EYfkavR8nW4Tb+AMkbfUFqmE6
l1bOI5o4FvEUbOxAsdC+1L0WfjsSucAenYQOCKROjVhNp7gjADGwnzjioMzE6+Rt7+uSiercFr8+
eLCingkxy1YZer0WRNGBczb7hAlKiPK9+eMVt2mzMLpSfDNqr4LxdogSSZc0Rw+XcntNriR05Xo0
twKPx1IQXCbR2pless7PF1Cu+lgrJwRyqYriSX/lsR7m/8EuLwF0rr7hcGYnqnkbo4mSsXVUFAhO
+ANepXuGKr/OtlZVEyfw2X1p19lRSNPGkjgDbgznYk+uecd8JCZ/mkpj9AJ6zxKTuKfOTzXQ31eY
D0gu6lTOxYoN7dgGsaySyfbbxEh+lOiN1ic/RSgZFWV+YV2uU7xjiEV+CqG/eYd6zJwWcvXKGQhZ
qz+jwEeA+bFCFJgJDoVkJVM/iY6f3HqTB0a08lkPUhoklLZrgyU6sxefocZkI52FHRwsfDZcHZ/3
XfWNmunoL7WlILbHFFQuODLHjFYzZ8+ybZbKyYzoi8bJddQPL1DcEY+x+qn15mgL8MsGlXhWvNbG
xBYUXobh6oHalubKohxQ3eWQjLgmtk8Y9vAzzzHSX3q7Aqfm/JBaRhq+9m3wJGSYqMAi6C3EvAMk
sWIr5AE6EiuvaTIaPwApUOZEsyjcYfOu4Doi1NJ9lFRLvNCprJlbvMWoSP4320HP3cKvosGbAu8O
i7pwMu2a/b/kLFT9rPFNAWvrs3HjsI7yi24XADNTLpaOJM2lpf4dAzBLYa8+V/gphyQBhHs0e6be
KuxpL6Krn6eDO/ZnWLXOLwZFGEwwnLIE3b0R1DY8YNExUbSDQ6VNTzewMSdtbPa3BCzK5cRi9bQh
gcfpvD9NSrJpKCCc9dqkdcFw1xDK8GOvMW5fWqv8Nrrj9Xx+tihhGTtrbWgQKKAUU4SOt5cFqbRq
2o1Bcws9HnkFAH/7RdxSdl882iRzIucLt2s7dZ2pA4GEl9Rs9TEoA9wi5cfGhdu40ueYjr8CCpZt
Dr/IjU2+MEYJ0qNzvu0SUQMbW058x3Y1ddiZjqpcJA==
`pragma protect end_protected
