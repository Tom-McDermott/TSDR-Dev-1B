// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
QFGBVVeCtcybYS+nEsO3BIYfdPpk+NhI+pgOapSh1Z+7R+KkiQgSesIeDWFbSvqC/dkej2t609Fr
Qg0xc5vBex4qlC45HB1zp78GZGiEiB7747MRkVe9NDdKmdKvsUnTHAwSlj+crWbug8blVoQqh3UO
9AnqzpkQn0xsJX2mBEz62T4c3+2p89qL+AZw+goWXlS29COzws4P5ClGMtSGDdXb7GRv0B1lAzwB
9fXIbl56aY9QnlJmFbcJtLy5akh6uXoO1DAEzzaIRY9LVuWLO9ZhCr8G+v8vc+hYpNYTWFNQ5X3d
UPfy5soxR7RlvjALu7GdQrXJh8Uh506Lg2Lhqg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5088)
4Z+1wgtCegrzx+jf7XOFOMjjVO7ZwPRrUrV9UM/UW3MTKPSypuAlQlLBy5cRKEcGQ0iDhFsR0Bgk
7Rnadnr4m86Q9BbiY5F4migjAhQx8xJaHllmBfY1BS8LPhmVCUviyFWpvWY+hr4WUTzPOkA+BTWj
KiWRRJf4iYWGkA+Z4TrF9wObaWW9sMJJULPPHCas9iNIFhiU/oltzbBfuKRSME6bYj1wTLHPb4xI
4fbKKoRcRHFpL2/Xied9oWlZOPp6b1TWr+fSLb7wAh3elQvqcSekDpPxTAnV+s7fDRKyQpOoUMsa
6oVEwohW3xn91ZmQvXnwObSrIy5goxm6O3HFtafo2Ffe5CXBeqHhB+zkD77P7mTmCKWTh4+GWVOC
gmOGlG04shN6xbfa7GwBxcET/Sj+yisXzPpc1gCp4uibE/W9yYOQLBddem9Y3UFr3mokOmnDUWrp
ouWvLwk94RE3TslnRFFhJJwyrp0L8+PNheKbmvohXYTPHuM4fRdumiRMMazkKiWt7HEeNGLu3nCo
TIeEaOdWvLFeQd2KkhVJMi4UCodDHBqHU4Se0F6LV0wB/7TKcKLioK1bL6E4ZqPMJvRPwfCC5MrG
zJQq8QdKDsBNSl6QTxvEC+PA6dSeS+hIVyF7TOyd+JJTs08nmTWVSVOsNYJ6s+Fs4SYnFTK944/Q
JLswozlKVl+ztp1w8jMnsqSUb/cEP1kdGAxL72vIV4jvb80h6njSwmNy+el5b2gPsIyABQEKa6od
7T2AGwHM5hqIuJo7jpUShwjMfAlvt7hohBDOO2GmVzApERxqMpIOqOkOotHp6mIklzfPeJbFVswh
Kmt2fXj/Wfw0ZnKku6F/6qjhd2Edv/dQUL7rpFs54Hg1TEKnCnYPuUii6SC7UFA3C3tcwUj/bwWf
ONjNjYU1dB3UiruoReXHMjNyxbfDXvS1Sj8pBPqyZtj80FH9+CpfSRUGOmoWycpU+XiujLdwPdKr
TG2S+fE8Yf8miFo8nB1aDH3xYi6K20vpUn49x558e7VSaFX5dCfSO5KenXpPBtkCwx2JyWb1uV/n
qp7QqbvhLZwbpDZ1IAQlOM5E6XoFhWIgkxhzY58X4g4NQkj8NnhUkgLfCwOvKZgk9azmeaHIULyp
dySEUQ+mIqaFiqB5r6b1ggeaFli1gQ43MvOPt179PINhmhIQNPmD0iLHVwjDbIC3g1gPeAx4WsXY
yyQyBlT/ggUDE0Pq0Wm0X9Nnoxn4nN+icAdDgbAIXxcmNdFpA9XHYLRvfhdtlkPxWkU+qi0Vil4B
RRqhKBw3c34PraVe2tPNIk2ABGKjxZiZNAhjxWNc45KqPwAS+4n2QNiWs0XWcyzXw3RZVVei/pEl
+wVApxNvm3y/x4+UGN4ckNmfW7GShud+F7IoUzj9cv9MZtYxHNjYKu236moiw6ZMZCobPJGtWStG
VDMUOUDRTOU2KtVSsJ0D1MJUIhk6sKPaeftevTaotydAOJix+Z6c2oDgQQAd+wyWdg674orhZ7Lo
E9Ywk7VrI4b22i47vNNoJN0MK2kjNcfCP5zSRCt+EMw94PxfebGtkb2CCXFx/6jLi6Coa1WXb2kl
a2Vw208rnSQMLIh31MzOC/yKoX4pDl1SGGZ5Uyrzb91EDVjMoQxOkiuq4SNR3Z1cfYfLgYKHj9PN
ATC2silaSN232Rsiai7Ny2gaPnxL8gHBlHrUU3aj7YPnFGzd8tqh8bBSOoJx2TM3jtwyZ34L6KS4
7rs/oYG8BbgvPBbdJcgect0cezq4YS7u4Eu/rvkkW1N4trtzIH8Zy9PxOsygZQVADNYMKiPwItgH
qXUaj5rkeuC+pZKJ33Eeylk0e1/ZZpRvI46Jpbbz2rxrJ70Pb15A7ei3p85yTU8/p1cqJr5TX6sj
Z/TgJBjIPwZsK+xMRVG5ZcHYY5NAZ0bH6IfUvY7htqJ+N9IJVYSb9jkkLYKHuiIAed0aIM1TwyFN
eZLnrF71J4Jefzb/ndnaMoDXMNQzz0a+n5kpHte7P5rPh6xZmD0tgBj2nKqASt97vL5KtbvMsdq7
LbChoBqH1VpsCJ29FYdf8qFdzki8Z1XtivMu0sUbQHMwVSRKIt5oiJfC3V/lesvwFM0OW/iHoDtW
+VX/OBdt3yIbbbCUjD0XX7jKxBYZ0uF18enykrwMHJ0BhMt8+sEiCafoHy9FaEo1lbHNZltijJA/
Aa6a+dbrXM/5hkq7FPpxkA+GPFtEP+ZDMKX85Q/0JpNGw4Lo4J05DqtdFMVpNr8iYjVNyFfOexio
RsEq2m9R5yIt5FdVOP9V7Mnw6fQE56Znn70KdkVvjV/vehPpNDre2b14XV0J5MlNkxLYfjhciL0q
i0AA3otzewEcwtJ/zmVZClQd/UWKpJM0keAzxY3uHNb/y/cUqD0RCsyq72sQaYK5S7cbnd1AQHkh
4b9qm1Xne5ebNGMojzCo2R5VQIokpjuVI0EgB9oRoodxlCTPwQUAlTSEF9HSV10hhSYxVLS9SKUg
if5CISgCm4HLEbHAhug9tgZfQKDrDu131Of3mL5Ep8cKVqn3O8gk+qbgOftSK9n96JZT+UhfIPn8
9s6Jwo0fM2G9qrbVhp9F4nCaQNC+jwkB9cBitArmU6hgeA9/SCo8AMg8sqVUqhNMt8Fk0g+O/qaM
3bCM6AfxCX2mLJflwS1O24iYsm0X3fMoWTTCSOciJ3x0yRNlXHZXJ8KvggwYsIFJImb6cLZWdjbK
pmYvrGS/KewX8qCtbyTvWhC+UXFwojcB3IQCyx+9n1ziakYsMmKE5vYOfNw+DAe8Ss2t3grbmiru
tUQ5n0BDS2fgWLo15j7iMEvMB4B/olBO2R9/3oinico/mK+zrNMudYJkx2uzNaFYgO4oaD7ubTlL
RzEM9VPEOPceAWEuwjngf9mPtayIcBSzIGHieIklxPV65z+1AdQ+MvgLaZCsAT70tiPbYa1zQhbO
5qUJVmY1shXnn1tcBywzTpJRl5GbUVO0S22WyqBv67KckmpYIGxe2bSmh9ykaoMR8ePWKtjcsJBg
qOlpzoCG2ySTcCkxYIO7Nwsqx2OYZrMM43FR66PThzUeKELntk0OkOOOuc/tHPCNjynEaqloPVDc
w8DB4g3U3Jeg/5+gVmFZ7wOK4iOQ+GziRelAA9bViJ6F8CWr29qpqnP4cniT3YdDLkP5TU/GHm4w
7boZZV4b9O5V/XI7vphWFMGiiU/lBYFlcHlRV7E8at5ZIqe4mVCTgAPOSscLDlWmvhN6SVOtJuzl
Rim96C+fuCNC+KaTDsr3QKJQD9Xhd/YL2Q1TpjNmNvc9e/DiAolCelnlwyiQpBDECQH0a7yEuXdV
/kwXJejavLyFzRAgI+w0L3woSl0+O3NQYbVkB8utf2JyWWFKm509fbYuGbb5OiDNpFpa7R/2+tyL
T/0oSkacDhWfU2P+1HMDxTU18YaYUhtzeI0oOCCgmTitoIIRAAha2fBPSTAHzmt97rQM3DL2J/p4
riB4Hl9UJiimclDCcMiCNODIODfgkjTneEagPz0shWgoISa07ifRmM/7ngyKt0atERTdKvsWqSgK
DmhJjVZoXrbuMKvRvnE8hLrsnnIoKE63laAQ0H4ZWIqV91t7Wesb1eI3bL+5BQeCnjoe2GBBSfYV
/HGUwqYNHS0AhzFoOKtWRV/t8tveVY+twVSE7kiu0zDbOGTwTcOqGcA9i0Gi8Kxkp9VX3Gn72IMI
SNqWq+XyapTEvtAIab11i1m7BXCWLKzAhmgCNF7VIgv4+UmjAwIXthvbHdQKO6mp1VyRldVBkQeE
tiMZlHG2ZKIKd6Vwo0nu9yE8ZMnQZStA8qphJ0K+SlQBPtcp2Vt6AxmTCoDceEK0EU3kzCQuCLZX
JNJwY7gkVgImEmUy3q/WgDh9Q3wHjHZQ2D9zxcUvtYVN6s1FDJfGkB2HPjdW0tqvQj7EUgUihPwL
OvBF6utWsV7LiSjwyzvgtH0AIDRHhhQKxhJ+9Mdk29oipkg7Jim+DA4Xs55NwTt4SlJxOA6pPWZW
sI8gSCUsPCidAsLILZHJt4am8XsDwj/uU+F0u3IiHF+VDwlRGhA7F0miF+CEiAnUv1J6tKcz0Qoq
a4ZkXYgpJS8rH8Bin8Hpwcwla7UaCJ3uxtRAvfwhBuiXUNBQuN1M2Lq5lOQfcBuYVoHqutiHoCMw
8oQUydg3wTa8eczdHCy0UarR/I0NLoT4X3t8QWBj+ir4XvPE+ghqqEK3ih9PdFueZ6+ygOE4uGVV
RfB9RwAfjsJPRhBkAJoYdBDDo9IDE9TTnZjjyVeSRHsyyDNBfpn9ZnTSKhDaiuPqL0qU7c40JD5E
IlTbpEnC5aZV6wCZ1TPhYB9272l1CEmV31dk3+wa2t4H+a3e4DQshMhNKliJ5bN+OdNzhlbfMVHT
Kc0bPs7dvGyhUYMR0x1zm2puYJNZIvkPz6hid1ozAifves+anPkwIO7mfOjhXbngQc3lAaN9MDr3
EMflmu25mka8itFR56GMAPRx1pi6H9aebPA9Arf+GWfIIF8PHFIps5ckVSLndJO1PBFo2Rqzw8b3
4i0x3EQsDPGnkQKds2TZB9MAXVoP4giML1tsBnMVzrQwEaVUt6UGWPgXsA3EBhTc+dIZFTd687IK
x9ZbCv+e9gcKPOhpiRFU2EqUW6NyWSN+W0GxXOI/aftP49OwgoK+2Hxl8u7P9CnOddjEK9N3vGPS
Y+OysAYoVetB93vFyup0WQ2iIyezXYCcH8DvmukRM6NIZ6JzHprKyLa3JJBrgUjf8sUJI2lw2Lhg
8hJNry5xYrr2SsFsYBq1xTIPLTDX0Wj3QWSn659lMOa8jFNu0NkQyMxozs29HWkX2e8/gIEsORCt
cc3IQ/qIfu0e9s0xkPvPYYalhwTDiVqX+0ot6+rzxdFgJHBf6YhNTR8Xy9VX5OxMrv87yAAzer3J
EO/E+Zb/SGmV2+HIe06mIJ2oSsexQozHywOUosPiuWGFfnoHtq5yHX67LO2pMUrJgaM0/8SDcao+
WwiFYgG6g+OnlQt2U4ETYighnh3y7daaP6jZjG+2j1I/1JBqIpFq1S6X8HN/RFEiZ0Nl2xtU+MQb
FKE28pJvJ9wX31tB34fKNm5wwSkF+nGbJI6QzI/Y/APo2fLdv6HOQW6PCvZtAi9qFUTs4Ng+BrLi
ss6icri4sCK8KLV+I7hLyqQpWO69I5YjuriPi44L0G6XjuKBrjzUWaCyrEyObRetjDDtI8jTKj41
3mkaYhM+cZxS/V/6OMQpwZOmYC13bWsQsaslaicByRkIolGzV8/miSFWuxz/jNdvZl+j6z2TJDoB
79G6FhFCidEpP9z2Krxi1BPsTeQMlvPtEDlbu9rWdPpMFK3KcSLQc1VghlgMmAt1AISUGQLMb6ag
8HwUz/oyP1TBtgXde+dRsjAAURv5O//V1osxLn0q/yJ1eQFhX/t3uMu09HrlxA+FS0JpykYO87eC
AGuM+U85zWB4Ra+ogENWLkCtvFvccK1jbuHyVSrF0lrHviS3fh6duxVEzdPzUyEPeq6Wf9ePl3sV
7PsxvW4dJn7j5/lLFuSbO/CKit9tbdF1yxZdkv4wk/UkbnKxZeVmIfkaYJHzQMBMNa552OLJKBmG
rtCZYJar+/Qcanrf29B3GxjW3GvtgjNC/SHqSt+e16iC6CSlHkdOPfZjnq00v2+Mod9f/ZpnrgU9
WDiYYQ9DEMJu6NQFJ1YW8QHYU0uiaZYlPCAlkdLbjnfiPuFmN9WMm+nQYzVPKZGfVa01w/qk8OK/
iKqtqU3AgGLPgiv15J4iQKCPohkV57otejcOl40nUNfp/bE0G7GyFI3ZB9ylccdRBcVplGgW5yn8
Y7dtjwEMBRxyvCtmJsXHNUp5JchFIoQCo+NQGdaObTZ93PUwWv+UYe+S27k4ttevRTBPndUSEBLH
V84o+x2l8w9Rgt8qiwparyRUtIYeKBzXpYFnQe/eFu10+OQQzeFv9CRWdjIdr0EIdEDMobBuNL4z
t6uqCVTOAJyOPPMuRcDzvK6E+3AgUwQa9zM44mKugAruiqPmJj8RktjK3Cc0czxIv2ExWm9+iIxc
WX9ihA9ptlUBXG67OQHn9SNmkYNIu7w7nhxE96U9DTLa++oUvI+jEnWsyhoiegLf5eNIRzViTMc0
syMBhaPJetnEodE85GTgf/ziGBqIFBno2NjGf/4QN3X87w8P1cdCMalcJmZGdCahTV+6F4PK+LBN
wkmq7dpYK6ToPZQkKvRscR0e5jYBFUIBK3BmJnSVzw3pNHfFydUmy1TuvMHymcLfrfiQ3VyybeI3
1KYpVPHcwuPChUuWY0fozuf70jXgmbxLWxfH7miC2wyhWf6HQT2kLRoTMr/DIvuTRLm33DOCBN3L
B/JbbYIiNv1KVNUbJfUnKCRQ6I77GZymZGCX5DlZx07W9SYTPpHZmAzMcqDMFYY8nHPBXMXF2/dI
DtVGK56UBTBqmqK1dqtGJR7hicUL6ZUXySntHsaykx12z45JNWVvVoQluyagXgySHDH5+2tbr6Kv
o9zCeWLEn6qUVRBtSuMNF4YVIePQaqaUWXvbDeO68FPd/lgx+C5Hv2Qgb/Yqg0df3xz4QHdI+2oh
xa7kszkKYigROM/i6DVCRIXx5heMZ1+GWLcQmtb3W12Gl4m2KoXO6J08pBOh2zixy1v03d7bU2Ck
c4zJbzHaOvngO9S2TLhv66ITwKXNFPiHk9dZN34Ri7FpyQPcwl6bIAqwRCqffH1DQ8KSJ+rm3v1L
w59rndyubyVUoNcrD0tv
`pragma protect end_protected
