//__ACDS_USER_COMMENT__ (C) 2001-2020 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
//__ACDS_USER_COMMENT__ ACDS 20.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H=W_M;JH4EB%9+F42JM(3=+RA6T"'UG9/3%;U#5L:$C;P#BV'Z"4 G0  
H#)D!US1.^PQ6F'6$\L+5S"/=DUULVZX$OZ<DXV^(!*%^0)\P#/OF<P  
HD#CMCLZD905I745I.R)*B0\3G7\0PTFY"<8G?21.(N33.=,08FA'RP  
H)F5ZQ9'!IF=H<'%=@I%#;L\M_+&_K.DM^-8PVWNX4BC %K:PE!#*J   
HPK-1W+]2)#3'O[S1-#"@M-?N87O$22Z^Z7XAC2=T=DVS3#__<-"3-P  
`pragma protect encoding=(enctype="uuencode",bytes=11472       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@SS%)F^WKV*K;'"\1_>TIEHH?]3"H@^9%@^\@4;R>*O4 
@P*S;\R4< _\(KT J;#>/X8](=*N#."FG' ),$TPDFO< 
@0T5Z(>2^FK3N+I/*U,(K'9Z^GC$#W7CM-5!65O%')?0 
@.K!.*-;I[+/7X-479T2!\^ J*!-$D+<KLYW2>?-:-PT 
@7+__0!Z/"Z=,:)AUKOEV?VO P9<4OKUZ2XZ_%=,PPL  
@K[2V2L$2R&,0L" .XU"# ('+-4;,^F$(+*Q8(L<8=?\ 
@B-\F$0BR)  BX9W,V,#FLNM[&O+T??2%V&6;/+9\2ZH 
@>JBES,+OFF'4:6_M4/F&)_)J'RBKGNR-+4F_29*X\A8 
@_1?E% =&@>YW&RSI-U^KEO!BEOM-F#QTR^X,/N%'AS\ 
@J\9T (VX)'>\C&1>>AX_#XA >IG=*]TQ1]$Y)HV"<,X 
@'WMAZV/@D=F:6VW/H6/&X:-I&/B]BI6+TE7PI7V(AS( 
@[X.[K\5%EJ15L*.C\K<)CS8<+Q^41CU8I=:\J&,RCE( 
@U4QO!',P[(E/&^Z<*L+K$36WQ"=Y#1&ASS=%)3AI$AL 
@+[Y(J"X201SN0^KH6*6RH,<*6$ ?,G+#A)U;ZQK_,=P 
@Y T;7?0G<E1^*.Y\%1RNCEX>"1C7S0"41@7:H$C2<!0 
@NU$2^PZ[MXX!C,'/8!J^@_U)S]!K<RWGAW(5[T#Z/S4 
@O'2>094XOA3,Y.K=E^V+3$Q"'R(:YQ0X@[@Z%\')!H  
@$DS95Z7,*K?_5[F"3IHG821Q'O\<AFB9.&\<F&^-.50 
@LR*_=%,_5RBT:K=""):"=7U4/-?8E-6Y& SY)RIHDY0 
@213VN78'@A:V+4:H,,G3I#B1I.VIQ/?;[EOJ6 0$RW$ 
@&+=X'IK$MCKA &7P\5_R8EZF*,KOR8?'@JW]IA70M6L 
@>9.=%LO%^TOHTR.D>LG^"(S.+3P*R)D!TTN%A@DQ46, 
@P27>\:[/DB@W,0]5V1<C2^!3>S98';21SJ1_@K&I4QP 
@.:\JZE5S&C+;)Z3=_<R82Q+@LNPF.#-G,UZCK6>W&+0 
@[)_$-E/QT =F3&79]VSD/G\CV.+TA0+A-;""+.CE"J4 
@:V6_,1QC CSIASGZ$[9B4LI'>/>4?):9"0=$%0JE?YX 
@HN9W8):*2,[R'J;WJ,Q _I%RO2L3)C5%$T1ZQPP59Q  
@!]* 1J$7FGWLQ5Z7FZ0[0]B8%I">/463]F?? /I&.=L 
@/SB9\2X.R@N3*-PRK.7.^4QQB8)C_&7@<G9+:E>JD8L 
@\, D:#K.C1N187YY*;A/'Y.X%UO2&K2D&S>0T)+ WW4 
@V\RAW36U'6R4DTSH@?]@A@ZK#$R0J$QWHNCU=$N%P=, 
@%E"[B6O[&(1R8MM\US&E#$C9ILKDS]4'/39,WO<^VX\ 
@4#C"9'!Y3M7#O*&M=_U)MZ#+)M8VDAF_=0.SQI>3T\L 
@ .(QG>WO]..UQ8%LPP5?#/&])S*^^U*W+)Z0#(DLJ^  
@M>-5+S4G(Z<;EOI2Q6EZ):& UTW&EZ-?6P(0P"HUFLX 
@5HS2@V%+KF;?54Q?(>)I!>4[&)'="C%INDM2A4Q[C4$ 
@DE:7EF'@96(\-!'!6.A*.*F5JTN8A5DL%%Q :QP=[(T 
@%V5=V?G\_U2PI_F83B@P,&5$_?0$<Q^\<_&=3Z(>J6( 
@<!FP5>-?<TDK^)>5?&TLZ"9]H9VW:M-!GJC#NM'YK*4 
@T6<]-6.]V]!!8UQ-TX&O=424%<=/">G 8WNZDTF?Q"4 
@LJ"3]HS>13]+9&N>:YSHU+4D"4P;2CVFTISLC2SW/30 
@^;N 09WIASFA',UZ+W3G8]@TY4X=X 7T1(<=TIWM0.H 
@$N-%5%RT;@WNQCFSH,Z?91=^F[IT-:XUPLUQXTR080$ 
@A'.[-FXY.ZW1R/6#!=@TKY;H LOS*NI(QNE)<QU-6JX 
@U1@R$\NA1ETH"@$#*6BB"2!]S-I4("RDNB(\5>W5AK\ 
@;U+28!T@S"TBRLO%=U 'M1ZU<ZXRO H;X,".<00":X< 
@%BWSQ@=BYF!%@&BLS@E"N3<!CCNZ*90]6('21CC<JOH 
@L #=:&0@WM!)_*@?$-5%&[X>'%%PA,_0D%CTZ8<4DS\ 
@K8/NHE[9=),X;< 23<^]FS-5? MU'3F"!]$%T+1B*08 
@@NS?B@3RQ6"Z6,I]#;B8[(9-%&_H(^=%DM[UX42.*U0 
@#&H<Z((E65)11#*TZ;^V!5@)#5W8S_3FMX,?3W!=R^X 
@0N,?&AAJ9YE2!,J;N\\ PU8RBJ!DRF['7DXR#T-+PD< 
@N1;RN?0Q1AMZEB*HNVKU=3&@^R# O)1,1PQ^]SJFQ6$ 
@G39$76'<',(! -^:EU  ER<BDSND!13!,F8!7UU%QV\ 
@*:*K_T>7R6D54F(EB!&/DCX$GVL>?;$#VW%#LM$0<Q  
@3=PT7SGI=B?"63WQW'&8:L<A$4A"V+.BQFQ95KT,H D 
@ %]\)@C2FK;14+58I]4#(&1GF T2!)H%AO\3DZ<%.,P 
@H"3XQ7CFTKH*%GA+_V\J,W<_WR,#V%"9X8 D@=<7A0D 
@Q3KGGXNB[[.#-*6!"YX)X8)'^HZ$79U4NV=@!OBRR\L 
@Y#HFHA_="F?U0 GNMH /CV_8KMP8%K,#*G$XI01S.(P 
@ML))(DRN^%$QEJD26H8;X/I#B1?BB!;@H/ 'B?-V794 
@QHH:6O] TG:%/O5N+LB62WC*3>-(,)V]Y*H&AFPR)$8 
@-<S2#JINEC'M77T7>2+MF>I)C%W]_KG##@0(7_P7+@( 
@H*S>\N9("'A]?O<S7;(\)-)ZO97#Z L?11A?D/]<8F( 
@#XLW'?#]P!%*1SFDZ%I5Q@RH*O B#M7M& 0NTS>,"0@ 
@U>WUBKU5TAA4'7Z6/K!LF_1I TD%A'Q<WZR5WU5K+48 
@=LU&N+;H8PO'(X(:/ME>)T162/MA:(3UKDV&8DU#!F0 
@$[L^'"R[E<;]J9<ANN]\-ZDBLT56\0[1N6&-EVV#/4T 
@89L,S*G@A]2!AO&D!D#8F&D3?\6.5MS@ETVUIVQH@'< 
@LV+R"\&:JVJSZ4[$>VP-"<B_7//L\B%"CV_^Z.Y])>$ 
@WBQ;\8 >"5?ZY$H7XP000'=<3>GL^F0;\!".!99]4OL 
@Z2^3XA)/@[,AXWKF%"4HZ6#=^$LL")'G MTF*7DUKOP 
@_[A$8Q66-T69H%T<;?]3IVS!HN@V%5S:?2@A=J@ P%H 
@"W\9FC/Z?&Z\0*>/ ,62?:IRNO,X)W(%H->VMR]IY^T 
@=V]0W%[>\T(ZA^86:=./QXJ5)!(E@(J=GI6@PG&9_2  
@DPG)UX, 3ZCHV;NM<SD1UT4(J%EE]YX^-RC30U.97>T 
@3[QSO_WFQK/X\0S@:IV55%+5\=46&EEL,W&4>;=-;*H 
@S]RG-IW;/=9$>C/^_XNK37\('1UP1J#QT=AJ3-3KO;X 
@D5>_[-K@/&'=!0,@NP0-,-'ZZA=M);PZE<:2V69[MC< 
@24^DB+PS5+AI$V A$H*[JR=?"\0\/V\LWA(9+^Y/3^H 
@C1*"7I9+6(.#\;,*4[U9A!6[8!5*EZ\T=PV$<-L!\7, 
@?U^9;[,TZ<@@%IBN-8&@)EGS6,]?ABTQT<,B7YL?J9L 
@"5W+$,V!4VHI3KMAV!0KW@2X"*2,#@GFVJF.VNVPA_$ 
@DJ8P39OB. P& -@L+L*=W\9.LSKBLD%,EU"K_-3)V6T 
@WBD<(3)MP8GP (+91(M5!(#:=]04]H!_#K V"6RI74< 
@_])U%?K=&FU.PL4>E.;[I#@3#5Q-L6_!-1@E2Z[0E0, 
@]J + U%H_57\HZRM'<GRQ[?3/BGGM00J!@LA]P+Q'FD 
@20Q7A-.]0I#9&!35Z3A7/E7QT)TC=I!DCSQ!8-\+,I8 
@_H7 %ZKC[<^@TA;94/'/#D>>JO$P\F!+3$Q)[;[>##4 
@X\8ZN90EM^:R5GKZ!(4FTDD38$><M]OZH=,6GS!G3<8 
@LK.H&*YZ@"YLA,%$H=GW0Q"A3!G)"9TRZFE&*5!MDM( 
@P*4QO*'-3M#N@-6#6%+TB$H2572W]88Q%RP.FF-S#XT 
@WE,\N&5D6FSP2!4]!H1#!*G+[5V,&)\HBHGQW6EF7J8 
@S,;(S?BID-_P52Y_(E3T#9%G=-WR"8^7)9)P%%AZA 0 
@K/AA<,]"U45NTO(N\/E$0!SCRTR>2YMMJW] #S^*5TL 
@ -YQF@R>D-NX-3]IE\.L:L*4*:UKUB\]UEA,#ITJO#, 
@IT0)^72;*:?XSVX=5V8F[S_T&B-L$%QM)<D# K#9A7H 
@[:R;+5[/H3:"/$68[?H)X.P9OL^J^][0I8<1QZ( H,< 
@=O7OAB.X%:)QL3BDQE7H SD#Y@+.!\+0M@B%F' M=U4 
@0BC#&^WPL2UT2HIMUWQ9\P! R9(TZ>T8?K[)+#V!F]@ 
@:YO=D_)UD*R%K37$KI-)Q>U9L>G4WNG!0@PTU1-"#64 
@C7T4B-MLBCBJU]'6&D-EXZ!HZWWA)MH>,T:0H$X,M@( 
@W9!H%JMK\=LN/+&X,/(7X-.CD='LL>C^;3E:3_;9#>\ 
@1]W#?^*>#E(MLB=H["ML=]+R-D4VI@AD9' 9W::[5=8 
@%?7WUG&9'>8UM=B6; 0@VXO:9=M,$4CUZ[:Q^S:FH>H 
@6=-YZ$L3_3L.$FDFU\BF*LLYCPKH@:N&5BN"7!KPW0L 
@CK\OKBZ5\@C.:S\-84V-Y^""/;2UW)0J[WJS6*NH%I< 
@IS4#SU2+;6I58 B[M 1 =V:1JS-A&R^NA.\^:AX9AIH 
@056U%4DNR(A=NT%).)1T+=%(OZ.Z)UG3"'Q><<0H 0( 
@#E@Q2G$ZOX"N</-5-N6$S&J79$U:!,_^&%EW('_)@!X 
@H>I!\9E\-]_E)::XF C5@I#VH_XM8(J=[.:B]<2I?'4 
@6V[U[R7-=DO_E9AJK\LP/6K,\@WH&.5.1. NR;*\GP@ 
@="?%DN6/;,\DT45%-NX\NS?L13Q?MF"Y-X\!PY"L]S( 
@ E']8-T1U8X>@$.;B"?QV\[1.F\9.O\8CN)\TABY(D( 
@. 8ND M6,\+6C1!Y["#DJD3PH4;.G]R[A-5M%GB037, 
@E3PZ8)VRT\_H2*H"1PYQ?6++;99Y=GFVG%#&I '+)8H 
@;.R"[@WE]<SUKT/;[T>65H+A20!>F@X%6(8E4+A-V<P 
@^*F[[_'RT0O1NVL) %0$3J0JAZ#D1U8(0BLP<(KRU@H 
@S*2.^O -GV!P)]^A-I]OZZ(M\\2XV$ ,F\8(FA$8PF( 
@)]R='AN,#[?J"@!*$"XC?VB4P)G7ZOK(O\I?X'%=P0< 
@/6K)HI=AZC-S&)3=%R:7_2!= (AK4]0>L,PZ_&6)\8< 
@A9P$3CYPIN19HL-4B+..U"K@;B5.V[$P_S$,/W.Q97L 
@BN*Y(D&F_'W6:=",PQTBFL-D[^J]EQK7HBUSJK\N)U@ 
@BQ0FO,>OD5P="R=3\T+NNK8/^G"0>#B,C NP38K I0, 
@#BN/].G.Q7@@DB"(( G)H,U(DF?P=,2= =EED!BYPBL 
@3I5(> / H$ K0\>%C [W"<00R('CF^,.&GQC1'>F,;T 
@,<MH6/D6C'TBI/;&"PM>%K0!IC'EKE=J\/:LVU]( F( 
@U";2H"I&@$QPI5,L:5!GXXM:F^B8_G;U1Y;U[<T'-?4 
@HU7=Z RD#*+2794M:$V4P'D:ID<9 &X8I,.G_8X<8R@ 
@OSA=/EME)[O$2Y(?N6)8L7[(4DR4A><P*L/$;+;7$70 
@'B^R6*H;,HSR1I$H;M-O[$,96CME!)%V/[#'AP76L8P 
@NA1\A=HN6_"."UAB?3DEC3HT[0WQYU68J=A-C"Y5F5D 
@1J7J87W^D&9 )2YG%T_4]'T\MUW,"T*$BR'G3@-G-&  
@U-<Z>#4_,,07MP093U\C>3A^0!R<\6MXX*)VT4,B>8$ 
@96>KWC%YC.8I-=U4>1Y(%7H?^[H#Q10<S(VP:3OC;>$ 
@(.C6?&=GC&25N$"*T<WBJTK%6N$T&SODC=!_-5A.TF\ 
@EO2+GH%!S*:_^5'&D1(1Y#[9*8C3RK8_/XYTP 4]#+$ 
@V$:UL 2P[U+[]4N<&8]833?SK<SYF/+*ZM$"P&UHR8T 
@U1H5L14CR(PX8-W,KR\HKA8<1DM?M'6ER5#\G,'(-&T 
@B=7,)V_[<@[-D9R?><'=[@NHN#>S1.[\Y\_0MBUJ$&P 
@*D-!P"H>GKR$C-6]T< )P)L-<T1[-L=%1E\6GUPF[\T 
@;@Q3U-"A\!N.;\)CZBSR@S*VZ&5C+^!^,#59]W*>YNX 
@&0*\%K';#+<M8RO-$T039JL&0R]"YYHFIEUM$B0LNI\ 
@3AZO4P4YB7*:S#G6#V$#<LL4,'T40/^%<BR9:#<MQQ$ 
@#;+%W1[9;##965B+-#QH_.+HR?_J?JMM3*QK&3?D[WT 
@8C;>=@6JUD$W# G!Q4\]=+,Q?FCUZ_J9-8DLHI@@:V4 
@+?]U'/+E$!9C0YW[HLAVS""W8B06+V-4E!0Y (U5[S0 
@G!._9]W=1 AL[3@"% .V4Z80Q+=<[EZRD6CRM!6X(+< 
@8$*',,'&%^4A";DEM7F[+5/Q-7FI;(RTRYYVSRJ5\C< 
@D @KFCI@E9SR^N:T2'CG: &*43HC=Z>/.)<@::G8.+  
@N+_L3E>GU3[;HI72N2N)+&*UYR+=L>8- #3@%:8QXX4 
@X7=)6:]+M[$*!0'!K I!5Q[WZS_6\6,UB+!^["JK33X 
@INW@(P(%5@;7\@ 'S>>)L__VHL4QFY2=F:U*9V8N^Z$ 
@>%FQ[U^(P+TM_+DNG>5YBT3<HV'3=$GWP;1N=-$\07\ 
@HD7/1MDA%C)#K>LY*JAG<A9_L(ONJ8-Y$3!OGU)!4?8 
@84-L7*/FJ,$N%27:Q3*(XK]0NN3G:* O!!TAJ$+$49L 
@Z4(>V,@-;+27%WK3_?,[.GBW'(""*0CJ?#X(2I:Q&PT 
@^;I L%"5!(,1G\Y]UK=2G5DGJ^PTQPZ)AH\.>=[?K^P 
@92!'0%&SHCT9!N/L%B$;\Y7'&NW$$'2'?:M*40$HBC( 
@ 7W2F%HEK-03,XZ?G7(J. F(,84 ^A_X9N7;?F7PF34 
@' Q_S"2C[&?ZY@3A):>LY3FHZ'RB_7JL1[D]^A Z'P0 
@_-^CRJ6Q]-M2C:_ZT!JP16<K[>3NY'@T:6E>8Y6(4:X 
@%@< X985T'/ZC2=O?IU[\M'P OY'=T-2!4L(\_R\DF4 
@J7)VD6B6#Y9&VAYC[L=7QG<;]JGV<L1LXW)H3Z\Y64< 
@Y$!:+@4TL?*#]3/A5>].&:%I4PO>&MN3/U3@!N.;MD4 
@E\@X>KN/BZ-",7_X  MDDZ13,O2G-0L@RB/QL#"XD+( 
@(YVK80WJ7WB#;5).-<U]YSH3-!1K?8.7R?P9-*%%LG@ 
@85;5YMDIK;&[BSRA2.E?MU5I#UT$'EO<M$,U C7$Y^D 
@4[F=:)O(L.\O^M_&6(\^1-P0'T<(Q-)R(,IT;GQ&:10 
@"@>%>YT\PON%?OE.%MH:HJIGFWUZ2D-[04.J%.;_E$T 
@J2?&67TX(P2L 07BI2:/+JP!QLRZL)TD&)C.H$>K#+\ 
@TN4$%A:<,UYQ/[>72K5XHOL_@WYV&P),1)'VH[X!X?P 
@@*&TW0BQC.4]XN.\3Z'UWV>]J)5G-&)0Z"GXJD+MX8X 
@47[(13=]B/V'@"N1<D4P;"M%=@EWISZG]:QP<MR!*\8 
@0R1V!$5T%>9!(U6'BWH)[OXHXC!N85,K>,0^=3*;_D( 
@?^,C^Q69CIK4#LLJX<#X<[&R172.X;0]=YJFI_;*Y H 
@,FTZUY+O<#RPC>J[2&1OBXZP8-P+OPZDRD6&M-;I/;X 
@B42L6 7F>X6-7T."4>T8H@#<:DX+( 9 1ZGAO__"1!@ 
@*1O'W)+_SXA0^B;&*4__Q3.Y3EOF3ER[46='&RKIH"\ 
@,OZ"5^Q[@,N*R%??V!(F0E()Z[9F(KYN/7ARNH$,D$L 
@?L/B-<<$1%KO^4Z&[ETX%E;X5*T3((:]&WD]H,4N\S  
@&:&ER_J08L'-C11(?Q&K4<$>:QKAC@(J-Z8ZMF,E/!  
@Q!6M9R%4> MHF/!;]DD9 /PN^$DOC]]H ;O^.ECQ62D 
@2F:G ]2+\!+[P](A%&+BVK@S\\]#Y=-/7>)-VJM<U:\ 
@>*Z8V3@42V)X/KA/$Z5%.HH6E0A<NH?>V+.51IJ1C8\ 
@*[S$Y#A")SH3 TWYZ[*F\5!>"!28)XI+2BGT'=HN1U( 
@QR+DT%I@@J5R E@"&%5MG)=^6(#U%X)\U5?EQ0GUG5  
@M6I<B/RUVL<[A:U0>"H'I6( X3TQ'[>01R"_L_/4RP8 
@3W>:<>Z1//Q/0P:&86^C4.4XFQS@^8@]0(A,\M#&W@0 
@5A$,A;Z*UL2C1'Q)@N0%F14X6F)0+!N:]Q= X]P5'<\ 
@)((N2U*I  8?=C(#\XB_T?I[8<&/2YZ+N? ZYX%RO\T 
@=A+ZYH2^Z$K2DDF&-R]ZZWVO!J$=JCC:.DL$=AA@:PX 
@2D.?SJ6IMNT@1)#L3;;D"]-6\8@LMZ3/*>ZKAW3U;>\ 
@R,&<"\2>'8U!I*;Q2[$3 N>FQM_[&G[S@KQ#!)D:PU4 
@EEZY90Q$%F*B#Z*+45$+,4/0:G5V],O+RX&SW4K5*\X 
@CL>69/F$2)FD6,X ^MD?> \\PT^>L-Z5O(N#"E]UQ\$ 
@WC#I<-,'%!,%,KL_E_@]6.SN[IX;O;$NM["!F=I9%9T 
@FS1;R+A[FIQGVU:FWTQ/$;]Q\ KL0O6(2H-@)J!3J7L 
@W53B3R0L&UOM*Z5>F4PQ;Q:E"+<UR63K4X N+XSI;/, 
@=W%AKBPLO"VT3K,[K;7#"ND"4IF^#]5@3/9!U*D<>N  
@I.9$Y^^DWU,77X :@Y<UO!PG6UERWDHKO#J/C\O?H@L 
@V@:%I[$U[WE;%T')_6%3K'\ MOK.8SS_+D)+KANH16X 
@"SKH@ /OE!0=I!4DSMA^&/#!.US[EHO4CS^_IFVM .H 
@K^&>%JQWKD9+A 'L'X)A0^Q>6ADX#0!PV * IN;HV)@ 
@KPQH^"'!P_L8=.]YX(>Q$ZWG^"FA/$T?+!<3:Y1=BB4 
@JX&F>?/.M[EG&%W*R +RR ,#?8!,FR=-WX9,K:W.O)D 
@NWE2@SUK/8%5NU18ELNK?%>3L+66#4AD!F&EF==[[=$ 
@0X+1/W/'Y&&B*C B$4"=UD^],SF,_J@-NO_&:G>RE$$ 
@'HN\>Z""U]NMXG*0:A42)Y;FAW\,^LG^_JIQX\B9UT, 
@$K"DNOX*##\^I;G+3'>#5F\;A>RFN7= F?G\AG:LU[T 
@/U:YE-1P_L*_Y^L7BN7(9RQ>N/.'!0I/$](P568W8G< 
@8RH:YIEUN&IO6\4EXG07-[[HZEC^$"U7DVROKU@8KB  
@YYK77*X]R->3*;-7"4V_F/W WY.#+\=4IIOD^QGP[]L 
@T#5XM?EAN\$$I:Q^S!+^QNUD@*5*7]9&29JYHH#2@:X 
@5;N5^*;9LF3-5(72- 9G(HJNZ.G<Q]9(MG.XJ3OC3FT 
@@FZHBYQ&C%"2>4.RCK&58<COKU2<Q^^V_>XPU+*9M(T 
@BH;YI<GZ-24Z2=OKMUY+MM';)>."K?K"[JAEECX&B38 
@Y 8E1CX><X^3-(DK!;JS4IB?4 9!4,ZUO"KF]_Y^%L8 
@*Y[H#9*4 /,C1U)J03='--F?DC?3_I(R!X#S(Y4%H0( 
@2!JQY0='COA>V1E6%J#C6T#LJ2_4EB-<W_''  K!)+D 
@FUZ4A4'>H_ A^+X/(5OGW+1R:/F,I+R0M-9WAO QOZ( 
@.P67W (U/ FB&;K!F[:\=WS.FPZ,X=P-AXJLTXV_?)H 
@95<(QLSVJWDXP5]H\OL6C;+ ;=^'E6L?$\G\=J<Z(W$ 
@AG1VBG-:7PQR1:S$.,^CG*',%J[NW5'M6<4AQY&ZV_0 
@_$5O3M#0./-+)P=D*HD&$,D9B1J!<G9L+WCR<TQ9P$D 
@A'NE(@XMXLHQU*WUN(B4ITWPZB&21R^#CF-\Y+GZJ54 
@<^+]<@:5_\D6R-;Q/MR*S=_X:0BGG8+^DJ6B@ZN#4$T 
@G-:"B#F@HA1PJU')B;H(#E..^M4!&0*+^?*7$0]EF%( 
@21&B#02YQ_8@I=&+^(2(\:J@N-IT#;R*8P3#HOJD/T4 
@G/M-@Q8X6:@0>U1';(*W8L!;S3\?.>WV[WEH#!9*/P4 
@ />\,F0>F1RIHY'M>1 J2O#@/\V@(.EX.,,MZ!C* DT 
@;"3YXQ PKM)[O8 KWEDR4,+O>.KO7/@R,*/ :B-$6=  
@P9< A 9K ;+&4B(>AO/O#HHG4^&- DQ,Y5=4#X-8QJ8 
@2G!@Q,YSSA0'DBD)_RUL!^;@K 7VIX[" 9N]E!19R^\ 
@?$?J=M>:,I=;7AMD8S*>P%.1V>C%2<I/57VR[Y;QF8H 
@:&O*>Q#;FS76!FAKLQ\KJV=C_( 1X.H;H=AT0S:VI(L 
@>YC F7+_-C08NJ9_,&L,W#FQ13 O])2],E&X:N-MY(( 
@-%%A#^4V?RFR"JXS%O5#9"ZO-UM7'X3ZACHMLH2-&+H 
@1E<&GM*SX:G?NDK@]6:[@+=%0M\U 98.$Y&6%K5IB*L 
@46X#>GU5N.W]/;FO+4#%-> B;*;"U$\I5=]IH>J)4"X 
@YM_RE 7"^&3,_,O4' 8E=?02_4O(E7OT1H85$^K1:M, 
@P;H69UAU8*[ZSM#ZD'5S5MO#=[6=2G9W9,X(F2D-048 
@<4+H$7YTE6"<SM!@<+@;YH1:CT!;#WE-!4[/%@VKQ/H 
@KP"AA%,"X:?MM!*H8(6%*B..= 7BOND"VS'#J1,%"G@ 
@^<VV!MT2[)"8)Q;-R 7K8Y&(Q'+G4"-I.$?.R>"[CX0 
@,!^$=VKPL_$NI![3]8H$S#V-8J7P]9,<K]D=8YMU9 X 
@N7GD$><G5B@$D$A_"5IH^Y-"G&0KV*"GT,(B +1D0GX 
@Z3ML[G4+6ED3#]/TK\YC>01.M2E]YWJV5>(O8KIK!P0 
@O4/T>(#'I$>KN<7>-RQ%L&RMR:#RCTHG!81+XKOP=3P 
@GYGA,S-H;,ZQO$SQ?0W^PL9R5)E=C-:P="D2!\^.OIL 
@0KM9-$1"RTJ,66-;EJ7M7O\_39&2,:XB?> K.0ID<7< 
@7YH<CB-&V[(ICAEISES=V65_$<4EP"^8&FQ0E?NTZ14 
@CE:$NV@+R#XEE3W'-CP4E2Z$![7'U"<4HLC8CZX)S4P 
@67RWLAPF)$6?M$YP!_UKQW<CC>B_/$6D/'^]T2Z5P*0 
@- ]H5 QFG[4U0&O9R>/X=Z@IJ<BKBF;,9K.NT(O):F\ 
@M\H'-(_^M3\+FEH T!RHB&K0!%8=O3G7!'B C>_)&Z0 
@8_D@E":%AY^EAI[X"57R=1*3;RNM-_<C-D\&$"P\M[, 
@3ADA-O7Y&><$P;E*X^7S*@+5:^^6I.4IL$34M;5T[%@ 
@D0X88V.GUGQ;VB9S2+TYR>[=ODL4J(,=+R WV7+C\?$ 
@G<&- 6H>BZPFDXR9;.U<R9R'A=* $#$JK@L>R!J%%AX 
@G"?JR+L>3.&[ZX,BA&5PCL6H.),V@TNUSR)2/QF1D1, 
@U5&4^^1Y22O11G.>.E<:T4&6:UQ #WATJ+-,"TL$8TH 
@8-*''$931]SLO/C2\ON4P"2OI-!_C@R=)![&,U0IR"\ 
@[\!@GWVX2Z!7!'U<8QEU,,(!B4[8+-%_;Y(17G@$/\L 
@EUN=/ZC&ION.(GP%;,&0&H>7'[B:!(K=+"ISE8*M3Z< 
@7M1B;XZR_C]/5*8S/]$%_8SCPYX[CK%D)@_*G5;.Q@@ 
@'FE%P<BCOW.D2<(AYUO=0K[;/FP?#F%"-)8-2Y*.#$T 
@>]U2_IX#[2F#9Z<VZH_AXFV2HI:ASY=2NZ>H&XM9I%8 
@IU;QO&FT$AH4)J80WM91(=:;&!]2^!V)"-8C^\4#QLD 
@2S)US4(26G99HYZ/"R !U6)N1K8&\2Q7]X7)[@AYZN  
@3L* 0@!BB].=Q#N"%JC%?[V9L')P9B72-:J!7F$ 2T8 
@BAQK^7GX^IC7,TB#CS:L]QHJITM*WD-P"%\>UL0+)=L 
@V>7W)?9'?3B4;QZDP)GM6N_+/SLN+PXFY:#B<=LBPCD 
@.HU=6+..9*RIHRND<FD%#HE1%V),T#D_%>RX+=1!70@ 
@WCWM\C8ZR\Q?9T5N2\.78([V.:Z5^FTP1Y/.^!O=J!P 
@@2^42\&G*0MO&0=$KJN84PZ$?KB1GXBBK-U$E(*?0SL 
@S<^K(26\$9;,['VI:-C^T\>Y)NBZ4$-WFLDDSN!.*M$ 
@Z@LPG^Z,FAQF/L)=M;S<\Y@/'C$V<".[8P+N__0%'!0 
@D!'&4Z-=GBY\XDDAC_&*M!,->WYH5K9-]3&EK<J/V$P 
@>U;98@A:S9DDLI[A(V41%N/K!+B5#II81O LG,L-7Y4 
@%=GEX\H0L_8[^[S[SYN6TAS1RV=,">EHQE7U(]Q6TV( 
@L^<6&521.CH;<F'J! !I3/'EH,J<7$PEP4O59$P<T \ 
@)[*OS=1<[CN@)G3VMXY,WR5+W4!5FCYRE:TT0>[98=\ 
@XCC4+IA\6\*JYH:P'EN'9+&,=2M8R:C1L.H<PK5L(NL 
@-QZ^<#@%F8U)#.?N(>1J")HPFOASU6MH1\"E$J,U-=$ 
@_H/P8/.F?E57K[B4SKG5I-G'#WU^/W-=LQ#B1UC=,<  
@N(OSYF' >):Q,95'#J;ZW^(&)FF@(%S/0=2>" Q'PV4 
@3*.BO]_Y:9ZXVR9!@C?!1$7X\'$=58^+B)@ON/MD\(H 
@I(2S;*+J22VPBP0#ST0>77_Z7I/(L;YW#(=4HZ\;ODX 
@FBH,91P8<CQM"Z-9A&Q!\U$4^/&+WAP/MDMLZN2L2$8 
@"BL\F;0F)K[I0/@$PSH,:@+9CW>PB;"7^)7[\.?W4%( 
@7E]>5\GKC&(=AR6[(]K$588L >=E)K/U"4D3VQL1/[  
@^;%XTQ8D;E98+5$-YDG4]_TK&2-B>[1"=ISFM9<:(FL 
@2N&KMK=$ -MLFL'PA@<T2M4UTH%OW*&/9EO]((LBZ^0 
@5WYDF=I80M:8;RQ5B3-YU(0B+C,LUB["@*64*.-+3J< 
@F6)$UK?"%M)J_19BP5]!-"ZE)+] ;G53="\99DJ':$H 
@S1FKR&F]3#,MDAES@ZFL*7MT)SKU($)J22]A8-;3N!  
@'FPDE?A5&9K<J_E;[BI[ECD:39 +V3QH!=Q>]2K!MN, 
@%M+-CH-,R:%%-8Y[9HYG'F4%;"U1^:?#.'"@U6PJM8< 
@-J@H;WM[M[!!V%O)-6%PWQR0;W6C5]V]DG0>^"#S"_< 
@+\\EL^"\?$W(-'Z1X2&8[);J:NQ"@;+PI@U^* =_5>@ 
@?_VKD T)G$QQ^%Y7":LDNC^N^S>S[ ACI:JCGBC<@;0 
@7A)U>HP#<+J&F4D,<UKF5UR4K#G:K)&OB2JZT*(=8LX 
@D0[#IG<+7;3C<./+7J5:M$L8K7KQG8;],P7[A-:B8JD 
@D1=3G+/NK:? J \6H*9EK:#(TEUI.A(-HI;JU.<LKRT 
@Z ,J%H]E>UR,_V_>A+X?Y/>CE1L0.XWPKK"\3__O )D 
@S$9O*]H71Z/A(PX#]XJ7KT 38#<#[H[02.R5P^X#B&D 
@-4[-# C1$5V:EP?UB=LSE@89MEV_D0SHT!FQRA.0OI, 
@83=FIT.1O]:^]I!SP]T/\<<0%AA#"KFA!JOY40T+ Q$ 
@?TQ$95GA(M35"I-"7VOAFFBNG'J*\^F=8I:.__,,NO< 
@W0$S80#RU = J0LJW*8%W.@G$O<^$_>OH=07%"JGLD, 
@ Z(C S5'(F(4&$A:RW\ET\.EC8S,=3GP&@'XH4/OY9D 
@JW>GQH:I!42&R$0X#;MI;K87F>_$%47Y,OK+1.#G8F4 
@LAWTR2$'"7?[X[K3^].RW,.^A%K;+4=/H.IFO7" *00 
@5R_!GC8\BDSW>?0QP?6D=.3[\!4<*(=?0(+,[/)DF   
@S44:]4WR/S7EKU-9H)10UD)Z''$@IEREH.+*Q;";.14 
@JH]9.^1KPXZJ%5%XTJ_>?$C9O9P"/?>K8X.>$5?O "H 
@"/AY:S5> TK7M];BJ "SWOM&P^_N:M^[:5W#FN..*88 
@PH%$6X8(?9NFB^ 2Z6MLI%.<6:./?MA@/2"H"2(4!D  
@MC&MZ?"8XVH+@4X");#DN3!..#[G?EM^;]?JYQB2V,, 
@@PM8F)W2FQ&&/&WB19@B+.OT@X-+5D>_K_V.(W'4 6T 
@2_F[4,2@*3"S(3V;M!K\A8"JR&#]5U@"A20\8SGD1ED 
@-'9YU010A0UDB19TS'08^%DPZ0ZG<QU^F6)FS$3I6Y< 
@O&6 JD,E:OC/.)6H>)>+IA0J+C&B0 ".RGM0 @@]K=  
@'>&Y#AR?=-=BS9%X&T"5YCJZ/$0JEK0"*K8B/[&7#LP 
@#R]5<G\_*S-/<?=T1MZ+Y!>$<<N'.I+:1<5\-\#(OOT 
@A.TOX4HODR&;--PR&*' L6U X @+W&V&_2:3*5W NCD 
@$J))8P(7(*H^)Z_P-,#6&+GX(E_@(C,#D?*P9!96P)< 
@'#5?;3FRMV+'P%K,[Q<*B.LV1M.UFZJ+3%IT52J_Q0$ 
@J3;!"D0GB6\4_WC%623JBO"(M*,U P*;_'?#GCQT^YH 
@0#3H,1AZRTF QYU2/$FMKF._Q(QF*[>]TN]E8/*J6"P 
@^1T";#;27>W0ODS_T,2SN1)+JK@7BW /[%W49NC-D.  
@Z%;?>(GM\D9S_A?&H]3HS<J6)^P!-/^FX<K7%)OY8(P 
@9QV=-BL\:LF.+!R=E1 #2WB7*K<WSDK\M&\U4$F2]K4 
@T#3W \9W(Y@K:&RL]ZX*LPY,IY-8WHY[CRRW^JB1Q.P 
@/>VC:73U.X8N<XOBUCN!H!X=\N4^,O!G1 #(X  88%< 
@\":_@_/EL@-ZY'G)<JBAQ4Z#',)$'=N!)N^H/T@.'MD 
@K'R36Z,PG1*YJ].!% 'TXR:^3W>/ET]EEFU*[XQL0 8 
@P*]N9'@3RJRVRH2<D(M=M>65(7IN#NBTHC+M 12S%C\ 
@FNJ5_M2]S7:1GY:LB=AH]*VQ>G?%;X[699?H79_A2Z8 
@MBQLW.(8?K(LTJ/&OMGW->RT!L<-[:<AF9WWR>2>.FH 
@[KNP+H'25RX8H4*SU;AQDN(424H5#71YP+J0 E#ESNL 
@%/[ 3%6TIYV4\V_>C*TD[NL(O8>PV)]K=EM;GT/B&I( 
@C ]MUVU+W;EF 3#P^@O[:_7T4^Z7+AE1F(DT[^.Z!>$ 
@Z0M5<G04B8R,7%MJY!F7+PHK"[]D^[3R:.]+QS#"G($ 
@CEB)9HY?80*=O. &-#J#&#--8W1C!1W@2.X0Y4?6:2$ 
@09M[&$N(_H=%-W#U@!8UTC&CX/;KA%_V61:G"YFF$:H 
@GD*1<T9-VP??5WU7^$.RUSAUUVC+"$1J0Q0,-Y&WF+< 
@S?:1#.'2I;Y&#R8'*Q;P2H[;UZ#2"/,>-_$=7[NH"_L 
@Z:N8(^?Y5N-[)Q7NIF@2#]&]K&EQMN;QB4;FXD]%Y,T 
@,!6GR*;%&L0"VU=8.IC$T&$1".YBS)];M3D[E]QG#L$ 
@UY90I[LY]3$VXYRZ'0*!,[*=LOQTSRSO_ZXB5J.U^", 
@03S1A1=(9)$H8Q28ZYW)$0B)OZ9.T#JVN:B]H1H8A1  
@:W/C^N]<$"\&;]Y@6YC=#YD1=&\UO>:_5^W[@YG  )P 
@%#HT]9;_=IZ%[F:!94":!?6UPP1$G<VH0L"WO>!0TF4 
@F+/ 0.*)@;5)UYPMYXX2?R>,^&285";Z4LZ*A\VS5R8 
@A7./?42Z*B,?*5-GJ5PFB!Q:8G K8_M9YQT"78R)%B@ 
@6R%'?^.X_/-*Z&VGZ;-@@T8^W+L.\VV=;BK:+@M5-,$ 
0-R,!DUW1LO72 1GGZK#$EP  
`pragma protect end_protected
