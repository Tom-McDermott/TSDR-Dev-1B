// q_sys.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module q_sys (
		output wire        altpll_shift_c0_clk,                         //                     altpll_shift_c0.clk
		output wire        altpll_shift_locked_conduit_export,          //         altpll_shift_locked_conduit.export
		input  wire        clock_bridge_0_in_clk_clk,                   //               clock_bridge_0_in_clk.clk
		output wire        enet_pll_c0_clk,                             //                         enet_pll_c0.clk
		output wire        enet_pll_c1_clk,                             //                         enet_pll_c1.clk
		output wire        enet_pll_c2_clk,                             //                         enet_pll_c2.clk
		output wire        enet_pll_c3_clk,                             //                         enet_pll_c3.clk
		output wire        enet_pll_c4_clk,                             //                         enet_pll_c4.clk
		output wire        enet_pll_locked_conduit_export,              //             enet_pll_locked_conduit.export
		output wire        eth_tse_mac_mdio_connection_mdc,             //         eth_tse_mac_mdio_connection.mdc
		input  wire        eth_tse_mac_mdio_connection_mdio_in,         //                                    .mdio_in
		output wire        eth_tse_mac_mdio_connection_mdio_out,        //                                    .mdio_out
		output wire        eth_tse_mac_mdio_connection_mdio_oen,        //                                    .mdio_oen
		input  wire [3:0]  eth_tse_mac_rgmii_connection_rgmii_in,       //        eth_tse_mac_rgmii_connection.rgmii_in
		output wire [3:0]  eth_tse_mac_rgmii_connection_rgmii_out,      //                                    .rgmii_out
		input  wire        eth_tse_mac_rgmii_connection_rx_control,     //                                    .rx_control
		output wire        eth_tse_mac_rgmii_connection_tx_control,     //                                    .tx_control
		input  wire        eth_tse_mac_status_connection_set_10,        //       eth_tse_mac_status_connection.set_10
		input  wire        eth_tse_mac_status_connection_set_1000,      //                                    .set_1000
		output wire        eth_tse_mac_status_connection_eth_mode,      //                                    .eth_mode
		output wire        eth_tse_mac_status_connection_ena_10,        //                                    .ena_10
		input  wire        eth_tse_pcs_mac_rx_clock_connection_clk,     // eth_tse_pcs_mac_rx_clock_connection.clk
		input  wire        eth_tse_pcs_mac_tx_clock_connection_clk,     // eth_tse_pcs_mac_tx_clock_connection.clk
		inout  wire [3:0]  ext_flash_flash_dataout_conduit_dataout,     //             ext_flash_flash_dataout.conduit_dataout
		output wire        ext_flash_flash_dclk_out_conduit_dclk_out,   //            ext_flash_flash_dclk_out.conduit_dclk_out
		output wire [0:0]  ext_flash_flash_ncs_conduit_ncs,             //                 ext_flash_flash_ncs.conduit_ncs
		output wire [3:0]  led_pio_external_connection_export,          //         led_pio_external_connection.export
		output wire        mem_if_ddr3_emif_0_status_local_init_done,   //           mem_if_ddr3_emif_0_status.local_init_done
		output wire        mem_if_ddr3_emif_0_status_local_cal_success, //                                    .local_cal_success
		output wire        mem_if_ddr3_emif_0_status_local_cal_fail,    //                                    .local_cal_fail
		input  wire        mem_resetn_in_reset_reset_n,                 //                 mem_resetn_in_reset.reset_n
		output wire [13:0] memory_mem_a,                                //                              memory.mem_a
		output wire [2:0]  memory_mem_ba,                               //                                    .mem_ba
		inout  wire [0:0]  memory_mem_ck,                               //                                    .mem_ck
		inout  wire [0:0]  memory_mem_ck_n,                             //                                    .mem_ck_n
		output wire [0:0]  memory_mem_cke,                              //                                    .mem_cke
		output wire [0:0]  memory_mem_cs_n,                             //                                    .mem_cs_n
		output wire [0:0]  memory_mem_dm,                               //                                    .mem_dm
		output wire [0:0]  memory_mem_ras_n,                            //                                    .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,                            //                                    .mem_cas_n
		output wire [0:0]  memory_mem_we_n,                             //                                    .mem_we_n
		output wire        memory_mem_reset_n,                          //                                    .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                               //                                    .mem_dq
		inout  wire [0:0]  memory_mem_dqs,                              //                                    .mem_dqs
		inout  wire [0:0]  memory_mem_dqs_n,                            //                                    .mem_dqs_n
		output wire [0:0]  memory_mem_odt,                              //                                    .mem_odt
		input  wire        reset_reset_n,                               //                               reset.reset_n
		input  wire        sys_clk_clk                                  //                             sys_clk.clk
	);

	wire         sgdma_tx_out_valid;                                          // sgdma_tx:out_valid -> eth_tse:ff_tx_wren
	wire  [31:0] sgdma_tx_out_data;                                           // sgdma_tx:out_data -> eth_tse:ff_tx_data
	wire         sgdma_tx_out_ready;                                          // eth_tse:ff_tx_rdy -> sgdma_tx:out_ready
	wire         sgdma_tx_out_startofpacket;                                  // sgdma_tx:out_startofpacket -> eth_tse:ff_tx_sop
	wire         sgdma_tx_out_endofpacket;                                    // sgdma_tx:out_endofpacket -> eth_tse:ff_tx_eop
	wire         sgdma_tx_out_error;                                          // sgdma_tx:out_error -> eth_tse:ff_tx_err
	wire   [1:0] sgdma_tx_out_empty;                                          // sgdma_tx:out_empty -> eth_tse:ff_tx_mod
	wire  [31:0] cpu_data_master_readdata;                                    // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                 // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                 // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [29:0] cpu_data_master_address;                                     // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                  // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                        // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                               // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                       // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                   // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                             // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                          // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [29:0] cpu_instruction_master_address;                              // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                 // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                        // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire  [31:0] sgdma_tx_m_read_readdata;                                    // mm_interconnect_0:sgdma_tx_m_read_readdata -> sgdma_tx:m_read_readdata
	wire         sgdma_tx_m_read_waitrequest;                                 // mm_interconnect_0:sgdma_tx_m_read_waitrequest -> sgdma_tx:m_read_waitrequest
	wire  [31:0] sgdma_tx_m_read_address;                                     // sgdma_tx:m_read_address -> mm_interconnect_0:sgdma_tx_m_read_address
	wire         sgdma_tx_m_read_read;                                        // sgdma_tx:m_read_read -> mm_interconnect_0:sgdma_tx_m_read_read
	wire         sgdma_tx_m_read_readdatavalid;                               // mm_interconnect_0:sgdma_tx_m_read_readdatavalid -> sgdma_tx:m_read_readdatavalid
	wire         sgdma_rx_m_write_waitrequest;                                // mm_interconnect_0:sgdma_rx_m_write_waitrequest -> sgdma_rx:m_write_waitrequest
	wire  [31:0] sgdma_rx_m_write_address;                                    // sgdma_rx:m_write_address -> mm_interconnect_0:sgdma_rx_m_write_address
	wire   [3:0] sgdma_rx_m_write_byteenable;                                 // sgdma_rx:m_write_byteenable -> mm_interconnect_0:sgdma_rx_m_write_byteenable
	wire         sgdma_rx_m_write_write;                                      // sgdma_rx:m_write_write -> mm_interconnect_0:sgdma_rx_m_write_write
	wire  [31:0] sgdma_rx_m_write_writedata;                                  // sgdma_rx:m_write_writedata -> mm_interconnect_0:sgdma_rx_m_write_writedata
	wire  [31:0] sgdma_rx_descriptor_read_readdata;                           // mm_interconnect_0:sgdma_rx_descriptor_read_readdata -> sgdma_rx:descriptor_read_readdata
	wire         sgdma_rx_descriptor_read_waitrequest;                        // mm_interconnect_0:sgdma_rx_descriptor_read_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	wire  [31:0] sgdma_rx_descriptor_read_address;                            // sgdma_rx:descriptor_read_address -> mm_interconnect_0:sgdma_rx_descriptor_read_address
	wire         sgdma_rx_descriptor_read_read;                               // sgdma_rx:descriptor_read_read -> mm_interconnect_0:sgdma_rx_descriptor_read_read
	wire         sgdma_rx_descriptor_read_readdatavalid;                      // mm_interconnect_0:sgdma_rx_descriptor_read_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	wire  [31:0] sgdma_tx_descriptor_read_readdata;                           // mm_interconnect_0:sgdma_tx_descriptor_read_readdata -> sgdma_tx:descriptor_read_readdata
	wire         sgdma_tx_descriptor_read_waitrequest;                        // mm_interconnect_0:sgdma_tx_descriptor_read_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	wire  [31:0] sgdma_tx_descriptor_read_address;                            // sgdma_tx:descriptor_read_address -> mm_interconnect_0:sgdma_tx_descriptor_read_address
	wire         sgdma_tx_descriptor_read_read;                               // sgdma_tx:descriptor_read_read -> mm_interconnect_0:sgdma_tx_descriptor_read_read
	wire         sgdma_tx_descriptor_read_readdatavalid;                      // mm_interconnect_0:sgdma_tx_descriptor_read_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	wire         sgdma_tx_descriptor_write_waitrequest;                       // mm_interconnect_0:sgdma_tx_descriptor_write_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	wire  [31:0] sgdma_tx_descriptor_write_address;                           // sgdma_tx:descriptor_write_address -> mm_interconnect_0:sgdma_tx_descriptor_write_address
	wire         sgdma_tx_descriptor_write_write;                             // sgdma_tx:descriptor_write_write -> mm_interconnect_0:sgdma_tx_descriptor_write_write
	wire  [31:0] sgdma_tx_descriptor_write_writedata;                         // sgdma_tx:descriptor_write_writedata -> mm_interconnect_0:sgdma_tx_descriptor_write_writedata
	wire         sgdma_rx_descriptor_write_waitrequest;                       // mm_interconnect_0:sgdma_rx_descriptor_write_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	wire  [31:0] sgdma_rx_descriptor_write_address;                           // sgdma_rx:descriptor_write_address -> mm_interconnect_0:sgdma_rx_descriptor_write_address
	wire         sgdma_rx_descriptor_write_write;                             // sgdma_rx:descriptor_write_write -> mm_interconnect_0:sgdma_rx_descriptor_write_write
	wire  [31:0] sgdma_rx_descriptor_write_writedata;                         // sgdma_rx:descriptor_write_writedata -> mm_interconnect_0:sgdma_rx_descriptor_write_writedata
	wire  [31:0] mm_interconnect_0_dual_boot_0_avalon_readdata;               // dual_boot_0:avmm_rcv_readdata -> mm_interconnect_0:dual_boot_0_avalon_readdata
	wire   [2:0] mm_interconnect_0_dual_boot_0_avalon_address;                // mm_interconnect_0:dual_boot_0_avalon_address -> dual_boot_0:avmm_rcv_address
	wire         mm_interconnect_0_dual_boot_0_avalon_read;                   // mm_interconnect_0:dual_boot_0_avalon_read -> dual_boot_0:avmm_rcv_read
	wire         mm_interconnect_0_dual_boot_0_avalon_write;                  // mm_interconnect_0:dual_boot_0_avalon_write -> dual_boot_0:avmm_rcv_write
	wire  [31:0] mm_interconnect_0_dual_boot_0_avalon_writedata;              // mm_interconnect_0:dual_boot_0_avalon_writedata -> dual_boot_0:avmm_rcv_writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;      // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;   // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_mem_if_ddr3_emif_0_avl_beginbursttransfer; // mm_interconnect_0:mem_if_ddr3_emif_0_avl_beginbursttransfer -> mem_if_ddr3_emif_0:avl_burstbegin
	wire  [31:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_readdata;           // mem_if_ddr3_emif_0:avl_rdata -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_readdata
	wire         mm_interconnect_0_mem_if_ddr3_emif_0_avl_waitrequest;        // mem_if_ddr3_emif_0:avl_ready -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_waitrequest
	wire  [24:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_address;            // mm_interconnect_0:mem_if_ddr3_emif_0_avl_address -> mem_if_ddr3_emif_0:avl_addr
	wire         mm_interconnect_0_mem_if_ddr3_emif_0_avl_read;               // mm_interconnect_0:mem_if_ddr3_emif_0_avl_read -> mem_if_ddr3_emif_0:avl_read_req
	wire   [3:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_byteenable;         // mm_interconnect_0:mem_if_ddr3_emif_0_avl_byteenable -> mem_if_ddr3_emif_0:avl_be
	wire         mm_interconnect_0_mem_if_ddr3_emif_0_avl_readdatavalid;      // mem_if_ddr3_emif_0:avl_rdata_valid -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_readdatavalid
	wire         mm_interconnect_0_mem_if_ddr3_emif_0_avl_write;              // mm_interconnect_0:mem_if_ddr3_emif_0_avl_write -> mem_if_ddr3_emif_0:avl_write_req
	wire  [31:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_writedata;          // mm_interconnect_0:mem_if_ddr3_emif_0_avl_writedata -> mem_if_ddr3_emif_0:avl_wdata
	wire   [2:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_burstcount;         // mm_interconnect_0:mem_if_ddr3_emif_0_avl_burstcount -> mem_if_ddr3_emif_0:avl_size
	wire         mem_if_ddr3_emif_0_afi_clk_clk;                              // mem_if_ddr3_emif_0:afi_clk -> [mm_interconnect_0:mem_if_ddr3_emif_0_afi_clk_clk, rst_controller_006:clk]
	wire  [31:0] mm_interconnect_0_ext_flash_avl_csr_readdata;                // ext_flash:avl_csr_rddata -> mm_interconnect_0:ext_flash_avl_csr_readdata
	wire         mm_interconnect_0_ext_flash_avl_csr_waitrequest;             // ext_flash:avl_csr_waitrequest -> mm_interconnect_0:ext_flash_avl_csr_waitrequest
	wire   [2:0] mm_interconnect_0_ext_flash_avl_csr_address;                 // mm_interconnect_0:ext_flash_avl_csr_address -> ext_flash:avl_csr_addr
	wire         mm_interconnect_0_ext_flash_avl_csr_read;                    // mm_interconnect_0:ext_flash_avl_csr_read -> ext_flash:avl_csr_read
	wire         mm_interconnect_0_ext_flash_avl_csr_readdatavalid;           // ext_flash:avl_csr_rddata_valid -> mm_interconnect_0:ext_flash_avl_csr_readdatavalid
	wire         mm_interconnect_0_ext_flash_avl_csr_write;                   // mm_interconnect_0:ext_flash_avl_csr_write -> ext_flash:avl_csr_write
	wire  [31:0] mm_interconnect_0_ext_flash_avl_csr_writedata;               // mm_interconnect_0:ext_flash_avl_csr_writedata -> ext_flash:avl_csr_wrdata
	wire  [31:0] mm_interconnect_0_ext_flash_avl_mem_readdata;                // ext_flash:avl_mem_rddata -> mm_interconnect_0:ext_flash_avl_mem_readdata
	wire         mm_interconnect_0_ext_flash_avl_mem_waitrequest;             // ext_flash:avl_mem_waitrequest -> mm_interconnect_0:ext_flash_avl_mem_waitrequest
	wire  [23:0] mm_interconnect_0_ext_flash_avl_mem_address;                 // mm_interconnect_0:ext_flash_avl_mem_address -> ext_flash:avl_mem_addr
	wire         mm_interconnect_0_ext_flash_avl_mem_read;                    // mm_interconnect_0:ext_flash_avl_mem_read -> ext_flash:avl_mem_read
	wire   [3:0] mm_interconnect_0_ext_flash_avl_mem_byteenable;              // mm_interconnect_0:ext_flash_avl_mem_byteenable -> ext_flash:avl_mem_byteenable
	wire         mm_interconnect_0_ext_flash_avl_mem_readdatavalid;           // ext_flash:avl_mem_rddata_valid -> mm_interconnect_0:ext_flash_avl_mem_readdatavalid
	wire         mm_interconnect_0_ext_flash_avl_mem_write;                   // mm_interconnect_0:ext_flash_avl_mem_write -> ext_flash:avl_mem_write
	wire  [31:0] mm_interconnect_0_ext_flash_avl_mem_writedata;               // mm_interconnect_0:ext_flash_avl_mem_writedata -> ext_flash:avl_mem_wrdata
	wire   [6:0] mm_interconnect_0_ext_flash_avl_mem_burstcount;              // mm_interconnect_0:ext_flash_avl_mem_burstcount -> ext_flash:avl_mem_burstcount
	wire  [31:0] mm_interconnect_0_eth_tse_control_port_readdata;             // eth_tse:reg_data_out -> mm_interconnect_0:eth_tse_control_port_readdata
	wire         mm_interconnect_0_eth_tse_control_port_waitrequest;          // eth_tse:reg_busy -> mm_interconnect_0:eth_tse_control_port_waitrequest
	wire   [7:0] mm_interconnect_0_eth_tse_control_port_address;              // mm_interconnect_0:eth_tse_control_port_address -> eth_tse:reg_addr
	wire         mm_interconnect_0_eth_tse_control_port_read;                 // mm_interconnect_0:eth_tse_control_port_read -> eth_tse:reg_rd
	wire         mm_interconnect_0_eth_tse_control_port_write;                // mm_interconnect_0:eth_tse_control_port_write -> eth_tse:reg_wr
	wire  [31:0] mm_interconnect_0_eth_tse_control_port_writedata;            // mm_interconnect_0:eth_tse_control_port_writedata -> eth_tse:reg_data_in
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;              // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;               // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_0_sgdma_tx_csr_chipselect;                   // mm_interconnect_0:sgdma_tx_csr_chipselect -> sgdma_tx:csr_chipselect
	wire  [31:0] mm_interconnect_0_sgdma_tx_csr_readdata;                     // sgdma_tx:csr_readdata -> mm_interconnect_0:sgdma_tx_csr_readdata
	wire   [3:0] mm_interconnect_0_sgdma_tx_csr_address;                      // mm_interconnect_0:sgdma_tx_csr_address -> sgdma_tx:csr_address
	wire         mm_interconnect_0_sgdma_tx_csr_read;                         // mm_interconnect_0:sgdma_tx_csr_read -> sgdma_tx:csr_read
	wire         mm_interconnect_0_sgdma_tx_csr_write;                        // mm_interconnect_0:sgdma_tx_csr_write -> sgdma_tx:csr_write
	wire  [31:0] mm_interconnect_0_sgdma_tx_csr_writedata;                    // mm_interconnect_0:sgdma_tx_csr_writedata -> sgdma_tx:csr_writedata
	wire         mm_interconnect_0_sgdma_rx_csr_chipselect;                   // mm_interconnect_0:sgdma_rx_csr_chipselect -> sgdma_rx:csr_chipselect
	wire  [31:0] mm_interconnect_0_sgdma_rx_csr_readdata;                     // sgdma_rx:csr_readdata -> mm_interconnect_0:sgdma_rx_csr_readdata
	wire   [3:0] mm_interconnect_0_sgdma_rx_csr_address;                      // mm_interconnect_0:sgdma_rx_csr_address -> sgdma_rx:csr_address
	wire         mm_interconnect_0_sgdma_rx_csr_read;                         // mm_interconnect_0:sgdma_rx_csr_read -> sgdma_rx:csr_read
	wire         mm_interconnect_0_sgdma_rx_csr_write;                        // mm_interconnect_0:sgdma_rx_csr_write -> sgdma_rx:csr_write
	wire  [31:0] mm_interconnect_0_sgdma_rx_csr_writedata;                    // mm_interconnect_0:sgdma_rx_csr_writedata -> sgdma_rx:csr_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;              // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;           // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;           // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;               // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                  // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;            // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                 // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;             // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_descriptor_memory_s1_chipselect;           // mm_interconnect_0:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	wire  [31:0] mm_interconnect_0_descriptor_memory_s1_readdata;             // descriptor_memory:readdata -> mm_interconnect_0:descriptor_memory_s1_readdata
	wire  [10:0] mm_interconnect_0_descriptor_memory_s1_address;              // mm_interconnect_0:descriptor_memory_s1_address -> descriptor_memory:address
	wire   [3:0] mm_interconnect_0_descriptor_memory_s1_byteenable;           // mm_interconnect_0:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	wire         mm_interconnect_0_descriptor_memory_s1_write;                // mm_interconnect_0:descriptor_memory_s1_write -> descriptor_memory:write
	wire  [31:0] mm_interconnect_0_descriptor_memory_s1_writedata;            // mm_interconnect_0:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	wire         mm_interconnect_0_descriptor_memory_s1_clken;                // mm_interconnect_0:descriptor_memory_s1_clken -> descriptor_memory:clken
	wire         mm_interconnect_0_sys_clk_timer_s1_chipselect;               // mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_readdata;                 // sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_timer_s1_address;                  // mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_0_sys_clk_timer_s1_write;                    // mm_interconnect_0:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_writedata;                // mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_0_onchip_ram_s1_chipselect;                  // mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_readdata;                    // onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	wire   [8:0] mm_interconnect_0_onchip_ram_s1_address;                     // mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	wire   [3:0] mm_interconnect_0_onchip_ram_s1_byteenable;                  // mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	wire         mm_interconnect_0_onchip_ram_s1_write;                       // mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_writedata;                   // mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	wire         mm_interconnect_0_onchip_ram_s1_clken;                       // mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	wire         mm_interconnect_0_led_pio_s1_chipselect;                     // mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	wire  [31:0] mm_interconnect_0_led_pio_s1_readdata;                       // led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_led_pio_s1_address;                        // mm_interconnect_0:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_0_led_pio_s1_write;                          // mm_interconnect_0:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_0_led_pio_s1_writedata;                      // mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	wire         irq_mapper_receiver0_irq;                                    // sgdma_rx:csr_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // sgdma_tx:csr_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver3_irq;                                    // jtag_uart:av_irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                    // sys_clk_timer:irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu_irq_irq;                                                 // irq_mapper:sender_irq -> cpu:irq
	wire         irq_mapper_receiver2_irq;                                    // irq_synchronizer:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                               // ext_flash:irq -> irq_synchronizer:receiver_irq
	wire         eth_tse_receive_valid;                                       // eth_tse:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire  [31:0] eth_tse_receive_data;                                        // eth_tse:ff_rx_data -> avalon_st_adapter:in_0_data
	wire         eth_tse_receive_ready;                                       // avalon_st_adapter:in_0_ready -> eth_tse:ff_rx_rdy
	wire         eth_tse_receive_startofpacket;                               // eth_tse:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire         eth_tse_receive_endofpacket;                                 // eth_tse:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire   [5:0] eth_tse_receive_error;                                       // eth_tse:rx_err -> avalon_st_adapter:in_0_error
	wire   [1:0] eth_tse_receive_empty;                                       // eth_tse:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                               // avalon_st_adapter:out_0_valid -> sgdma_rx:in_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                                // avalon_st_adapter:out_0_data -> sgdma_rx:in_data
	wire         avalon_st_adapter_out_0_ready;                               // sgdma_rx:in_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                       // avalon_st_adapter:out_0_startofpacket -> sgdma_rx:in_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                         // avalon_st_adapter:out_0_endofpacket -> sgdma_rx:in_endofpacket
	wire   [5:0] avalon_st_adapter_out_0_error;                               // avalon_st_adapter:out_0_error -> sgdma_rx:in_error
	wire   [1:0] avalon_st_adapter_out_0_empty;                               // avalon_st_adapter:out_0_empty -> sgdma_rx:in_empty
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [altpll_shift:reset, enet_pll:reset]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [cpu:reset_n, dual_boot_0:nreset, irq_mapper:reset, irq_synchronizer:sender_reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [avalon_st_adapter:in_rst_0_reset, descriptor_memory:reset, eth_tse:reset, jtag_uart:rst_n, led_pio:reset_n, mm_interconnect_0:sgdma_tx_reset_reset_bridge_in_reset_reset, onchip_ram:reset, rst_translator_001:in_reset, sgdma_rx:system_reset_n, sgdma_tx:system_reset_n, sys_clk_timer:reset_n, sysid:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                      // rst_controller_002:reset_req -> [descriptor_memory:reset_req, onchip_ram:reset_req, rst_translator_001:reset_req_in]
	wire         cpu_debug_reset_request_reset;                               // cpu:debug_reset_request -> [rst_controller_002:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in0, rst_controller_005:reset_in0, rst_controller_006:reset_in0]
	wire         rst_controller_003_reset_out_reset;                          // rst_controller_003:reset_out -> [ext_flash:reset_n, irq_synchronizer:receiver_reset, mm_interconnect_0:ext_flash_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_004_reset_out_reset;                          // rst_controller_004:reset_out -> mem_if_ddr3_emif_0:global_reset_n
	wire         rst_controller_005_reset_out_reset;                          // rst_controller_005:reset_out -> mem_if_ddr3_emif_0:soft_reset_n
	wire         rst_controller_006_reset_out_reset;                          // rst_controller_006:reset_out -> [mm_interconnect_0:mem_if_ddr3_emif_0_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mem_if_ddr3_emif_0_soft_reset_reset_bridge_in_reset_reset]

	q_sys_altpll_shift altpll_shift (
		.clk       (sys_clk_clk),                        //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),     // inclk_interface_reset.reset
		.read      (),                                   //             pll_slave.read
		.write     (),                                   //                      .write
		.address   (),                                   //                      .address
		.readdata  (),                                   //                      .readdata
		.writedata (),                                   //                      .writedata
		.c0        (altpll_shift_c0_clk),                //                    c0.clk
		.areset    (),                                   //        areset_conduit.export
		.c2        (),                                   //            c2_conduit.export
		.c1        (),                                   //            c1_conduit.export
		.locked    (altpll_shift_locked_conduit_export)  //        locked_conduit.export
	);

	q_sys_cpu cpu (
		.clk                                 (sys_clk_clk),                                       //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),               //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),            //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	q_sys_descriptor_memory descriptor_memory (
		.clk        (sys_clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_descriptor_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_descriptor_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_descriptor_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_descriptor_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_descriptor_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_descriptor_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_descriptor_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req)             //       .reset_req
	);

	altera_dual_boot #(
		.INTENDED_DEVICE_FAMILY ("MAX 10"),
		.CONFIG_CYCLE           (18),
		.RESET_TIMER_CYCLE      (26)
	) dual_boot_0 (
		.clk                (sys_clk_clk),                                    //    clk.clk
		.nreset             (~rst_controller_001_reset_out_reset),            // nreset.reset_n
		.avmm_rcv_address   (mm_interconnect_0_dual_boot_0_avalon_address),   // avalon.address
		.avmm_rcv_read      (mm_interconnect_0_dual_boot_0_avalon_read),      //       .read
		.avmm_rcv_writedata (mm_interconnect_0_dual_boot_0_avalon_writedata), //       .writedata
		.avmm_rcv_write     (mm_interconnect_0_dual_boot_0_avalon_write),     //       .write
		.avmm_rcv_readdata  (mm_interconnect_0_dual_boot_0_avalon_readdata)   //       .readdata
	);

	q_sys_enet_pll enet_pll (
		.clk       (sys_clk_clk),                    //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                               //             pll_slave.read
		.write     (),                               //                      .write
		.address   (),                               //                      .address
		.readdata  (),                               //                      .readdata
		.writedata (),                               //                      .writedata
		.c0        (enet_pll_c0_clk),                //                    c0.clk
		.c1        (enet_pll_c1_clk),                //                    c1.clk
		.c2        (enet_pll_c2_clk),                //                    c2.clk
		.c3        (enet_pll_c3_clk),                //                    c3.clk
		.c4        (enet_pll_c4_clk),                //                    c4.clk
		.locked    (enet_pll_locked_conduit_export)  //        locked_conduit.export
	);

	q_sys_eth_tse eth_tse (
		.clk           (sys_clk_clk),                                        // control_port_clock_connection.clk
		.reset         (rst_controller_002_reset_out_reset),                 //              reset_connection.reset
		.reg_addr      (mm_interconnect_0_eth_tse_control_port_address),     //                  control_port.address
		.reg_data_out  (mm_interconnect_0_eth_tse_control_port_readdata),    //                              .readdata
		.reg_rd        (mm_interconnect_0_eth_tse_control_port_read),        //                              .read
		.reg_data_in   (mm_interconnect_0_eth_tse_control_port_writedata),   //                              .writedata
		.reg_wr        (mm_interconnect_0_eth_tse_control_port_write),       //                              .write
		.reg_busy      (mm_interconnect_0_eth_tse_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (eth_tse_pcs_mac_tx_clock_connection_clk),            //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (eth_tse_pcs_mac_rx_clock_connection_clk),            //   pcs_mac_rx_clock_connection.clk
		.set_10        (eth_tse_mac_status_connection_set_10),               //         mac_status_connection.set_10
		.set_1000      (eth_tse_mac_status_connection_set_1000),             //                              .set_1000
		.eth_mode      (eth_tse_mac_status_connection_eth_mode),             //                              .eth_mode
		.ena_10        (eth_tse_mac_status_connection_ena_10),               //                              .ena_10
		.rgmii_in      (eth_tse_mac_rgmii_connection_rgmii_in),              //          mac_rgmii_connection.rgmii_in
		.rgmii_out     (eth_tse_mac_rgmii_connection_rgmii_out),             //                              .rgmii_out
		.rx_control    (eth_tse_mac_rgmii_connection_rx_control),            //                              .rx_control
		.tx_control    (eth_tse_mac_rgmii_connection_tx_control),            //                              .tx_control
		.ff_rx_clk     (sys_clk_clk),                                        //      receive_clock_connection.clk
		.ff_tx_clk     (sys_clk_clk),                                        //     transmit_clock_connection.clk
		.ff_rx_data    (eth_tse_receive_data),                               //                       receive.data
		.ff_rx_eop     (eth_tse_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (eth_tse_receive_error),                              //                              .error
		.ff_rx_mod     (eth_tse_receive_empty),                              //                              .empty
		.ff_rx_rdy     (eth_tse_receive_ready),                              //                              .ready
		.ff_rx_sop     (eth_tse_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (eth_tse_receive_valid),                              //                              .valid
		.ff_tx_data    (sgdma_tx_out_data),                                  //                      transmit.data
		.ff_tx_eop     (sgdma_tx_out_endofpacket),                           //                              .endofpacket
		.ff_tx_err     (sgdma_tx_out_error),                                 //                              .error
		.ff_tx_mod     (sgdma_tx_out_empty),                                 //                              .empty
		.ff_tx_rdy     (sgdma_tx_out_ready),                                 //                              .ready
		.ff_tx_sop     (sgdma_tx_out_startofpacket),                         //                              .startofpacket
		.ff_tx_wren    (sgdma_tx_out_valid),                                 //                              .valid
		.mdc           (eth_tse_mac_mdio_connection_mdc),                    //           mac_mdio_connection.mdc
		.mdio_in       (eth_tse_mac_mdio_connection_mdio_in),                //                              .mdio_in
		.mdio_out      (eth_tse_mac_mdio_connection_mdio_out),               //                              .mdio_out
		.mdio_oen      (eth_tse_mac_mdio_connection_mdio_oen),               //                              .mdio_oen
		.magic_wakeup  (),                                                   //           mac_misc_connection.magic_wakeup
		.magic_sleep_n (),                                                   //                              .magic_sleep_n
		.ff_tx_crc_fwd (),                                                   //                              .ff_tx_crc_fwd
		.ff_tx_septy   (),                                                   //                              .ff_tx_septy
		.tx_ff_uflow   (),                                                   //                              .tx_ff_uflow
		.ff_tx_a_full  (),                                                   //                              .ff_tx_a_full
		.ff_tx_a_empty (),                                                   //                              .ff_tx_a_empty
		.rx_err_stat   (),                                                   //                              .rx_err_stat
		.rx_frm_type   (),                                                   //                              .rx_frm_type
		.ff_rx_dsav    (),                                                   //                              .ff_rx_dsav
		.ff_rx_a_full  (),                                                   //                              .ff_rx_a_full
		.ff_rx_a_empty ()                                                    //                              .ff_rx_a_empty
	);

	generic_qspi_controller #(
		.DEVICE_FAMILY     ("MAX 10"),
		.CS_WIDTH          (1),
		.ADDR_WIDTH        (24),
		.ASI_WIDTH         (4),
		.ASMI_ADDR_WIDTH   (32),
		.ENABLE_4BYTE_ADDR (1),
		.IO_MODE           ("QUAD"),
		.CHIP_SELS         (1)
	) ext_flash (
		.clk                  (clock_bridge_0_in_clk_clk),                         //       clock_sink.clk
		.reset_n              (~rst_controller_003_reset_out_reset),               //            reset.reset_n
		.avl_csr_read         (mm_interconnect_0_ext_flash_avl_csr_read),          //          avl_csr.read
		.avl_csr_waitrequest  (mm_interconnect_0_ext_flash_avl_csr_waitrequest),   //                 .waitrequest
		.avl_csr_write        (mm_interconnect_0_ext_flash_avl_csr_write),         //                 .write
		.avl_csr_addr         (mm_interconnect_0_ext_flash_avl_csr_address),       //                 .address
		.avl_csr_wrdata       (mm_interconnect_0_ext_flash_avl_csr_writedata),     //                 .writedata
		.avl_csr_rddata       (mm_interconnect_0_ext_flash_avl_csr_readdata),      //                 .readdata
		.avl_csr_rddata_valid (mm_interconnect_0_ext_flash_avl_csr_readdatavalid), //                 .readdatavalid
		.avl_mem_write        (mm_interconnect_0_ext_flash_avl_mem_write),         //          avl_mem.write
		.avl_mem_burstcount   (mm_interconnect_0_ext_flash_avl_mem_burstcount),    //                 .burstcount
		.avl_mem_waitrequest  (mm_interconnect_0_ext_flash_avl_mem_waitrequest),   //                 .waitrequest
		.avl_mem_read         (mm_interconnect_0_ext_flash_avl_mem_read),          //                 .read
		.avl_mem_addr         (mm_interconnect_0_ext_flash_avl_mem_address),       //                 .address
		.avl_mem_wrdata       (mm_interconnect_0_ext_flash_avl_mem_writedata),     //                 .writedata
		.avl_mem_rddata       (mm_interconnect_0_ext_flash_avl_mem_readdata),      //                 .readdata
		.avl_mem_rddata_valid (mm_interconnect_0_ext_flash_avl_mem_readdatavalid), //                 .readdatavalid
		.avl_mem_byteenable   (mm_interconnect_0_ext_flash_avl_mem_byteenable),    //                 .byteenable
		.irq                  (irq_synchronizer_receiver_irq),                     // interrupt_sender.irq
		.flash_dataout        (ext_flash_flash_dataout_conduit_dataout),           //    flash_dataout.conduit_dataout
		.flash_dclk_out       (ext_flash_flash_dclk_out_conduit_dclk_out),         //   flash_dclk_out.conduit_dclk_out
		.flash_ncs            (ext_flash_flash_ncs_conduit_ncs)                    //        flash_ncs.conduit_ncs
	);

	q_sys_jtag_uart jtag_uart (
		.clk            (sys_clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                   //               irq.irq
	);

	q_sys_led_pio led_pio (
		.clk        (sys_clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_external_connection_export)       // external_connection.export
	);

	q_sys_mem_if_ddr3_emif_0 mem_if_ddr3_emif_0 (
		.pll_ref_clk        (sys_clk_clk),                                                 //      pll_ref_clk.clk
		.global_reset_n     (~rst_controller_004_reset_out_reset),                         //     global_reset.reset_n
		.soft_reset_n       (~rst_controller_005_reset_out_reset),                         //       soft_reset.reset_n
		.afi_clk            (mem_if_ddr3_emif_0_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk       (),                                                            //     afi_half_clk.clk
		.afi_reset_n        (),                                                            //        afi_reset.reset_n
		.afi_reset_export_n (),                                                            // afi_reset_export.reset_n
		.mem_a              (memory_mem_a),                                                //           memory.mem_a
		.mem_ba             (memory_mem_ba),                                               //                 .mem_ba
		.mem_ck             (memory_mem_ck),                                               //                 .mem_ck
		.mem_ck_n           (memory_mem_ck_n),                                             //                 .mem_ck_n
		.mem_cke            (memory_mem_cke),                                              //                 .mem_cke
		.mem_cs_n           (memory_mem_cs_n),                                             //                 .mem_cs_n
		.mem_dm             (memory_mem_dm),                                               //                 .mem_dm
		.mem_ras_n          (memory_mem_ras_n),                                            //                 .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),                                            //                 .mem_cas_n
		.mem_we_n           (memory_mem_we_n),                                             //                 .mem_we_n
		.mem_reset_n        (memory_mem_reset_n),                                          //                 .mem_reset_n
		.mem_dq             (memory_mem_dq),                                               //                 .mem_dq
		.mem_dqs            (memory_mem_dqs),                                              //                 .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),                                            //                 .mem_dqs_n
		.mem_odt            (memory_mem_odt),                                              //                 .mem_odt
		.avl_ready          (mm_interconnect_0_mem_if_ddr3_emif_0_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin     (mm_interconnect_0_mem_if_ddr3_emif_0_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr           (mm_interconnect_0_mem_if_ddr3_emif_0_avl_address),            //                 .address
		.avl_rdata_valid    (mm_interconnect_0_mem_if_ddr3_emif_0_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata          (mm_interconnect_0_mem_if_ddr3_emif_0_avl_readdata),           //                 .readdata
		.avl_wdata          (mm_interconnect_0_mem_if_ddr3_emif_0_avl_writedata),          //                 .writedata
		.avl_be             (mm_interconnect_0_mem_if_ddr3_emif_0_avl_byteenable),         //                 .byteenable
		.avl_read_req       (mm_interconnect_0_mem_if_ddr3_emif_0_avl_read),               //                 .read
		.avl_write_req      (mm_interconnect_0_mem_if_ddr3_emif_0_avl_write),              //                 .write
		.avl_size           (mm_interconnect_0_mem_if_ddr3_emif_0_avl_burstcount),         //                 .burstcount
		.local_init_done    (mem_if_ddr3_emif_0_status_local_init_done),                   //           status.local_init_done
		.local_cal_success  (mem_if_ddr3_emif_0_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail     (mem_if_ddr3_emif_0_status_local_cal_fail),                    //                 .local_cal_fail
		.pll_mem_clk        (),                                                            //      pll_sharing.pll_mem_clk
		.pll_write_clk      (),                                                            //                 .pll_write_clk
		.pll_locked         (),                                                            //                 .pll_locked
		.pll_capture0_clk   (),                                                            //                 .pll_capture0_clk
		.pll_capture1_clk   ()                                                             //                 .pll_capture1_clk
	);

	q_sys_onchip_ram onchip_ram (
		.clk        (sys_clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_onchip_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req)      //       .reset_req
	);

	q_sys_sgdma_rx sgdma_rx (
		.clk                           (sys_clk_clk),                               //              clk.clk
		.system_reset_n                (~rst_controller_002_reset_out_reset),       //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_rx_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_rx_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_rx_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_rx_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_rx_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_rx_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_rx_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_rx_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_rx_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_rx_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),                  //          csr_irq.irq
		.in_startofpacket              (avalon_st_adapter_out_0_startofpacket),     //               in.startofpacket
		.in_endofpacket                (avalon_st_adapter_out_0_endofpacket),       //                 .endofpacket
		.in_data                       (avalon_st_adapter_out_0_data),              //                 .data
		.in_valid                      (avalon_st_adapter_out_0_valid),             //                 .valid
		.in_ready                      (avalon_st_adapter_out_0_ready),             //                 .ready
		.in_empty                      (avalon_st_adapter_out_0_empty),             //                 .empty
		.in_error                      (avalon_st_adapter_out_0_error),             //                 .error
		.m_write_waitrequest           (sgdma_rx_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (sgdma_rx_m_write_address),                  //                 .address
		.m_write_write                 (sgdma_rx_m_write_write),                    //                 .write
		.m_write_writedata             (sgdma_rx_m_write_writedata),                //                 .writedata
		.m_write_byteenable            (sgdma_rx_m_write_byteenable)                //                 .byteenable
	);

	q_sys_sgdma_tx sgdma_tx (
		.clk                           (sys_clk_clk),                               //              clk.clk
		.system_reset_n                (~rst_controller_002_reset_out_reset),       //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_tx_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_tx_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_tx_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_tx_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_tx_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_tx_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_tx_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_tx_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_tx_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_tx_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver1_irq),                  //          csr_irq.irq
		.m_read_readdata               (sgdma_tx_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_tx_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_tx_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_tx_m_read_read),                      //                 .read
		.out_data                      (sgdma_tx_out_data),                         //              out.data
		.out_valid                     (sgdma_tx_out_valid),                        //                 .valid
		.out_ready                     (sgdma_tx_out_ready),                        //                 .ready
		.out_endofpacket               (sgdma_tx_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (sgdma_tx_out_startofpacket),                //                 .startofpacket
		.out_empty                     (sgdma_tx_out_empty),                        //                 .empty
		.out_error                     (sgdma_tx_out_error)                         //                 .error
	);

	q_sys_sys_clk_timer sys_clk_timer (
		.clk        (sys_clk_clk),                                   //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                       //   irq.irq
	);

	q_sys_sysid sysid (
		.clock    (sys_clk_clk),                                    //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	q_sys_mm_interconnect_0 mm_interconnect_0 (
		.clock_bridge_0_out_clk_clk                                          (clock_bridge_0_in_clk_clk),                                   //                                        clock_bridge_0_out_clk.clk
		.mem_if_ddr3_emif_0_afi_clk_clk                                      (mem_if_ddr3_emif_0_afi_clk_clk),                              //                                    mem_if_ddr3_emif_0_afi_clk.clk
		.sys_clk_clk_clk                                                     (sys_clk_clk),                                                 //                                                   sys_clk_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset                               (rst_controller_001_reset_out_reset),                          //                               cpu_reset_reset_bridge_in_reset.reset
		.ext_flash_reset_reset_bridge_in_reset_reset                         (rst_controller_003_reset_out_reset),                          //                         ext_flash_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_0_avl_translator_reset_reset_bridge_in_reset_reset (rst_controller_006_reset_out_reset),                          // mem_if_ddr3_emif_0_avl_translator_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_0_soft_reset_reset_bridge_in_reset_reset           (rst_controller_006_reset_out_reset),                          //           mem_if_ddr3_emif_0_soft_reset_reset_bridge_in_reset.reset
		.sgdma_tx_reset_reset_bridge_in_reset_reset                          (rst_controller_002_reset_out_reset),                          //                          sgdma_tx_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                             (cpu_data_master_address),                                     //                                               cpu_data_master.address
		.cpu_data_master_waitrequest                                         (cpu_data_master_waitrequest),                                 //                                                              .waitrequest
		.cpu_data_master_byteenable                                          (cpu_data_master_byteenable),                                  //                                                              .byteenable
		.cpu_data_master_read                                                (cpu_data_master_read),                                        //                                                              .read
		.cpu_data_master_readdata                                            (cpu_data_master_readdata),                                    //                                                              .readdata
		.cpu_data_master_readdatavalid                                       (cpu_data_master_readdatavalid),                               //                                                              .readdatavalid
		.cpu_data_master_write                                               (cpu_data_master_write),                                       //                                                              .write
		.cpu_data_master_writedata                                           (cpu_data_master_writedata),                                   //                                                              .writedata
		.cpu_data_master_debugaccess                                         (cpu_data_master_debugaccess),                                 //                                                              .debugaccess
		.cpu_instruction_master_address                                      (cpu_instruction_master_address),                              //                                        cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                                  (cpu_instruction_master_waitrequest),                          //                                                              .waitrequest
		.cpu_instruction_master_read                                         (cpu_instruction_master_read),                                 //                                                              .read
		.cpu_instruction_master_readdata                                     (cpu_instruction_master_readdata),                             //                                                              .readdata
		.cpu_instruction_master_readdatavalid                                (cpu_instruction_master_readdatavalid),                        //                                                              .readdatavalid
		.sgdma_rx_descriptor_read_address                                    (sgdma_rx_descriptor_read_address),                            //                                      sgdma_rx_descriptor_read.address
		.sgdma_rx_descriptor_read_waitrequest                                (sgdma_rx_descriptor_read_waitrequest),                        //                                                              .waitrequest
		.sgdma_rx_descriptor_read_read                                       (sgdma_rx_descriptor_read_read),                               //                                                              .read
		.sgdma_rx_descriptor_read_readdata                                   (sgdma_rx_descriptor_read_readdata),                           //                                                              .readdata
		.sgdma_rx_descriptor_read_readdatavalid                              (sgdma_rx_descriptor_read_readdatavalid),                      //                                                              .readdatavalid
		.sgdma_rx_descriptor_write_address                                   (sgdma_rx_descriptor_write_address),                           //                                     sgdma_rx_descriptor_write.address
		.sgdma_rx_descriptor_write_waitrequest                               (sgdma_rx_descriptor_write_waitrequest),                       //                                                              .waitrequest
		.sgdma_rx_descriptor_write_write                                     (sgdma_rx_descriptor_write_write),                             //                                                              .write
		.sgdma_rx_descriptor_write_writedata                                 (sgdma_rx_descriptor_write_writedata),                         //                                                              .writedata
		.sgdma_rx_m_write_address                                            (sgdma_rx_m_write_address),                                    //                                              sgdma_rx_m_write.address
		.sgdma_rx_m_write_waitrequest                                        (sgdma_rx_m_write_waitrequest),                                //                                                              .waitrequest
		.sgdma_rx_m_write_byteenable                                         (sgdma_rx_m_write_byteenable),                                 //                                                              .byteenable
		.sgdma_rx_m_write_write                                              (sgdma_rx_m_write_write),                                      //                                                              .write
		.sgdma_rx_m_write_writedata                                          (sgdma_rx_m_write_writedata),                                  //                                                              .writedata
		.sgdma_tx_descriptor_read_address                                    (sgdma_tx_descriptor_read_address),                            //                                      sgdma_tx_descriptor_read.address
		.sgdma_tx_descriptor_read_waitrequest                                (sgdma_tx_descriptor_read_waitrequest),                        //                                                              .waitrequest
		.sgdma_tx_descriptor_read_read                                       (sgdma_tx_descriptor_read_read),                               //                                                              .read
		.sgdma_tx_descriptor_read_readdata                                   (sgdma_tx_descriptor_read_readdata),                           //                                                              .readdata
		.sgdma_tx_descriptor_read_readdatavalid                              (sgdma_tx_descriptor_read_readdatavalid),                      //                                                              .readdatavalid
		.sgdma_tx_descriptor_write_address                                   (sgdma_tx_descriptor_write_address),                           //                                     sgdma_tx_descriptor_write.address
		.sgdma_tx_descriptor_write_waitrequest                               (sgdma_tx_descriptor_write_waitrequest),                       //                                                              .waitrequest
		.sgdma_tx_descriptor_write_write                                     (sgdma_tx_descriptor_write_write),                             //                                                              .write
		.sgdma_tx_descriptor_write_writedata                                 (sgdma_tx_descriptor_write_writedata),                         //                                                              .writedata
		.sgdma_tx_m_read_address                                             (sgdma_tx_m_read_address),                                     //                                               sgdma_tx_m_read.address
		.sgdma_tx_m_read_waitrequest                                         (sgdma_tx_m_read_waitrequest),                                 //                                                              .waitrequest
		.sgdma_tx_m_read_read                                                (sgdma_tx_m_read_read),                                        //                                                              .read
		.sgdma_tx_m_read_readdata                                            (sgdma_tx_m_read_readdata),                                    //                                                              .readdata
		.sgdma_tx_m_read_readdatavalid                                       (sgdma_tx_m_read_readdatavalid),                               //                                                              .readdatavalid
		.cpu_debug_mem_slave_address                                         (mm_interconnect_0_cpu_debug_mem_slave_address),               //                                           cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                           (mm_interconnect_0_cpu_debug_mem_slave_write),                 //                                                              .write
		.cpu_debug_mem_slave_read                                            (mm_interconnect_0_cpu_debug_mem_slave_read),                  //                                                              .read
		.cpu_debug_mem_slave_readdata                                        (mm_interconnect_0_cpu_debug_mem_slave_readdata),              //                                                              .readdata
		.cpu_debug_mem_slave_writedata                                       (mm_interconnect_0_cpu_debug_mem_slave_writedata),             //                                                              .writedata
		.cpu_debug_mem_slave_byteenable                                      (mm_interconnect_0_cpu_debug_mem_slave_byteenable),            //                                                              .byteenable
		.cpu_debug_mem_slave_waitrequest                                     (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),           //                                                              .waitrequest
		.cpu_debug_mem_slave_debugaccess                                     (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),           //                                                              .debugaccess
		.descriptor_memory_s1_address                                        (mm_interconnect_0_descriptor_memory_s1_address),              //                                          descriptor_memory_s1.address
		.descriptor_memory_s1_write                                          (mm_interconnect_0_descriptor_memory_s1_write),                //                                                              .write
		.descriptor_memory_s1_readdata                                       (mm_interconnect_0_descriptor_memory_s1_readdata),             //                                                              .readdata
		.descriptor_memory_s1_writedata                                      (mm_interconnect_0_descriptor_memory_s1_writedata),            //                                                              .writedata
		.descriptor_memory_s1_byteenable                                     (mm_interconnect_0_descriptor_memory_s1_byteenable),           //                                                              .byteenable
		.descriptor_memory_s1_chipselect                                     (mm_interconnect_0_descriptor_memory_s1_chipselect),           //                                                              .chipselect
		.descriptor_memory_s1_clken                                          (mm_interconnect_0_descriptor_memory_s1_clken),                //                                                              .clken
		.dual_boot_0_avalon_address                                          (mm_interconnect_0_dual_boot_0_avalon_address),                //                                            dual_boot_0_avalon.address
		.dual_boot_0_avalon_write                                            (mm_interconnect_0_dual_boot_0_avalon_write),                  //                                                              .write
		.dual_boot_0_avalon_read                                             (mm_interconnect_0_dual_boot_0_avalon_read),                   //                                                              .read
		.dual_boot_0_avalon_readdata                                         (mm_interconnect_0_dual_boot_0_avalon_readdata),               //                                                              .readdata
		.dual_boot_0_avalon_writedata                                        (mm_interconnect_0_dual_boot_0_avalon_writedata),              //                                                              .writedata
		.eth_tse_control_port_address                                        (mm_interconnect_0_eth_tse_control_port_address),              //                                          eth_tse_control_port.address
		.eth_tse_control_port_write                                          (mm_interconnect_0_eth_tse_control_port_write),                //                                                              .write
		.eth_tse_control_port_read                                           (mm_interconnect_0_eth_tse_control_port_read),                 //                                                              .read
		.eth_tse_control_port_readdata                                       (mm_interconnect_0_eth_tse_control_port_readdata),             //                                                              .readdata
		.eth_tse_control_port_writedata                                      (mm_interconnect_0_eth_tse_control_port_writedata),            //                                                              .writedata
		.eth_tse_control_port_waitrequest                                    (mm_interconnect_0_eth_tse_control_port_waitrequest),          //                                                              .waitrequest
		.ext_flash_avl_csr_address                                           (mm_interconnect_0_ext_flash_avl_csr_address),                 //                                             ext_flash_avl_csr.address
		.ext_flash_avl_csr_write                                             (mm_interconnect_0_ext_flash_avl_csr_write),                   //                                                              .write
		.ext_flash_avl_csr_read                                              (mm_interconnect_0_ext_flash_avl_csr_read),                    //                                                              .read
		.ext_flash_avl_csr_readdata                                          (mm_interconnect_0_ext_flash_avl_csr_readdata),                //                                                              .readdata
		.ext_flash_avl_csr_writedata                                         (mm_interconnect_0_ext_flash_avl_csr_writedata),               //                                                              .writedata
		.ext_flash_avl_csr_readdatavalid                                     (mm_interconnect_0_ext_flash_avl_csr_readdatavalid),           //                                                              .readdatavalid
		.ext_flash_avl_csr_waitrequest                                       (mm_interconnect_0_ext_flash_avl_csr_waitrequest),             //                                                              .waitrequest
		.ext_flash_avl_mem_address                                           (mm_interconnect_0_ext_flash_avl_mem_address),                 //                                             ext_flash_avl_mem.address
		.ext_flash_avl_mem_write                                             (mm_interconnect_0_ext_flash_avl_mem_write),                   //                                                              .write
		.ext_flash_avl_mem_read                                              (mm_interconnect_0_ext_flash_avl_mem_read),                    //                                                              .read
		.ext_flash_avl_mem_readdata                                          (mm_interconnect_0_ext_flash_avl_mem_readdata),                //                                                              .readdata
		.ext_flash_avl_mem_writedata                                         (mm_interconnect_0_ext_flash_avl_mem_writedata),               //                                                              .writedata
		.ext_flash_avl_mem_burstcount                                        (mm_interconnect_0_ext_flash_avl_mem_burstcount),              //                                                              .burstcount
		.ext_flash_avl_mem_byteenable                                        (mm_interconnect_0_ext_flash_avl_mem_byteenable),              //                                                              .byteenable
		.ext_flash_avl_mem_readdatavalid                                     (mm_interconnect_0_ext_flash_avl_mem_readdatavalid),           //                                                              .readdatavalid
		.ext_flash_avl_mem_waitrequest                                       (mm_interconnect_0_ext_flash_avl_mem_waitrequest),             //                                                              .waitrequest
		.jtag_uart_avalon_jtag_slave_address                                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),       //                                   jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),         //                                                              .write
		.jtag_uart_avalon_jtag_slave_read                                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),          //                                                              .read
		.jtag_uart_avalon_jtag_slave_readdata                                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),      //                                                              .readdata
		.jtag_uart_avalon_jtag_slave_writedata                               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),     //                                                              .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),   //                                                              .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),    //                                                              .chipselect
		.led_pio_s1_address                                                  (mm_interconnect_0_led_pio_s1_address),                        //                                                    led_pio_s1.address
		.led_pio_s1_write                                                    (mm_interconnect_0_led_pio_s1_write),                          //                                                              .write
		.led_pio_s1_readdata                                                 (mm_interconnect_0_led_pio_s1_readdata),                       //                                                              .readdata
		.led_pio_s1_writedata                                                (mm_interconnect_0_led_pio_s1_writedata),                      //                                                              .writedata
		.led_pio_s1_chipselect                                               (mm_interconnect_0_led_pio_s1_chipselect),                     //                                                              .chipselect
		.mem_if_ddr3_emif_0_avl_address                                      (mm_interconnect_0_mem_if_ddr3_emif_0_avl_address),            //                                        mem_if_ddr3_emif_0_avl.address
		.mem_if_ddr3_emif_0_avl_write                                        (mm_interconnect_0_mem_if_ddr3_emif_0_avl_write),              //                                                              .write
		.mem_if_ddr3_emif_0_avl_read                                         (mm_interconnect_0_mem_if_ddr3_emif_0_avl_read),               //                                                              .read
		.mem_if_ddr3_emif_0_avl_readdata                                     (mm_interconnect_0_mem_if_ddr3_emif_0_avl_readdata),           //                                                              .readdata
		.mem_if_ddr3_emif_0_avl_writedata                                    (mm_interconnect_0_mem_if_ddr3_emif_0_avl_writedata),          //                                                              .writedata
		.mem_if_ddr3_emif_0_avl_beginbursttransfer                           (mm_interconnect_0_mem_if_ddr3_emif_0_avl_beginbursttransfer), //                                                              .beginbursttransfer
		.mem_if_ddr3_emif_0_avl_burstcount                                   (mm_interconnect_0_mem_if_ddr3_emif_0_avl_burstcount),         //                                                              .burstcount
		.mem_if_ddr3_emif_0_avl_byteenable                                   (mm_interconnect_0_mem_if_ddr3_emif_0_avl_byteenable),         //                                                              .byteenable
		.mem_if_ddr3_emif_0_avl_readdatavalid                                (mm_interconnect_0_mem_if_ddr3_emif_0_avl_readdatavalid),      //                                                              .readdatavalid
		.mem_if_ddr3_emif_0_avl_waitrequest                                  (~mm_interconnect_0_mem_if_ddr3_emif_0_avl_waitrequest),       //                                                              .waitrequest
		.onchip_ram_s1_address                                               (mm_interconnect_0_onchip_ram_s1_address),                     //                                                 onchip_ram_s1.address
		.onchip_ram_s1_write                                                 (mm_interconnect_0_onchip_ram_s1_write),                       //                                                              .write
		.onchip_ram_s1_readdata                                              (mm_interconnect_0_onchip_ram_s1_readdata),                    //                                                              .readdata
		.onchip_ram_s1_writedata                                             (mm_interconnect_0_onchip_ram_s1_writedata),                   //                                                              .writedata
		.onchip_ram_s1_byteenable                                            (mm_interconnect_0_onchip_ram_s1_byteenable),                  //                                                              .byteenable
		.onchip_ram_s1_chipselect                                            (mm_interconnect_0_onchip_ram_s1_chipselect),                  //                                                              .chipselect
		.onchip_ram_s1_clken                                                 (mm_interconnect_0_onchip_ram_s1_clken),                       //                                                              .clken
		.sgdma_rx_csr_address                                                (mm_interconnect_0_sgdma_rx_csr_address),                      //                                                  sgdma_rx_csr.address
		.sgdma_rx_csr_write                                                  (mm_interconnect_0_sgdma_rx_csr_write),                        //                                                              .write
		.sgdma_rx_csr_read                                                   (mm_interconnect_0_sgdma_rx_csr_read),                         //                                                              .read
		.sgdma_rx_csr_readdata                                               (mm_interconnect_0_sgdma_rx_csr_readdata),                     //                                                              .readdata
		.sgdma_rx_csr_writedata                                              (mm_interconnect_0_sgdma_rx_csr_writedata),                    //                                                              .writedata
		.sgdma_rx_csr_chipselect                                             (mm_interconnect_0_sgdma_rx_csr_chipselect),                   //                                                              .chipselect
		.sgdma_tx_csr_address                                                (mm_interconnect_0_sgdma_tx_csr_address),                      //                                                  sgdma_tx_csr.address
		.sgdma_tx_csr_write                                                  (mm_interconnect_0_sgdma_tx_csr_write),                        //                                                              .write
		.sgdma_tx_csr_read                                                   (mm_interconnect_0_sgdma_tx_csr_read),                         //                                                              .read
		.sgdma_tx_csr_readdata                                               (mm_interconnect_0_sgdma_tx_csr_readdata),                     //                                                              .readdata
		.sgdma_tx_csr_writedata                                              (mm_interconnect_0_sgdma_tx_csr_writedata),                    //                                                              .writedata
		.sgdma_tx_csr_chipselect                                             (mm_interconnect_0_sgdma_tx_csr_chipselect),                   //                                                              .chipselect
		.sys_clk_timer_s1_address                                            (mm_interconnect_0_sys_clk_timer_s1_address),                  //                                              sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                                              (mm_interconnect_0_sys_clk_timer_s1_write),                    //                                                              .write
		.sys_clk_timer_s1_readdata                                           (mm_interconnect_0_sys_clk_timer_s1_readdata),                 //                                                              .readdata
		.sys_clk_timer_s1_writedata                                          (mm_interconnect_0_sys_clk_timer_s1_writedata),                //                                                              .writedata
		.sys_clk_timer_s1_chipselect                                         (mm_interconnect_0_sys_clk_timer_s1_chipselect),               //                                                              .chipselect
		.sysid_control_slave_address                                         (mm_interconnect_0_sysid_control_slave_address),               //                                           sysid_control_slave.address
		.sysid_control_slave_readdata                                        (mm_interconnect_0_sysid_control_slave_readdata)               //                                                              .readdata
	);

	q_sys_irq_mapper irq_mapper (
		.clk           (sys_clk_clk),                        //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (cpu_irq_irq)                         //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clock_bridge_0_in_clk_clk),          //       receiver_clk.clk
		.sender_clk     (sys_clk_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	q_sys_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (6),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (sys_clk_clk),                           // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_002_reset_out_reset),    // in_rst_0.reset
		.in_0_data           (eth_tse_receive_data),                  //     in_0.data
		.in_0_valid          (eth_tse_receive_valid),                 //         .valid
		.in_0_ready          (eth_tse_receive_ready),                 //         .ready
		.in_0_startofpacket  (eth_tse_receive_startofpacket),         //         .startofpacket
		.in_0_endofpacket    (eth_tse_receive_endofpacket),           //         .endofpacket
		.in_0_empty          (eth_tse_receive_empty),                 //         .empty
		.in_0_error          (eth_tse_receive_error),                 //         .error
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)          //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~mem_resetn_in_reset_reset_n),   // reset_in0.reset
		.clk            (sys_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (sys_clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),          // reset_in1.reset
		.clk            (sys_clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clock_bridge_0_in_clk_clk),          //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (cpu_debug_reset_request_reset),      // reset_in0.reset
		.reset_in1      (~mem_resetn_in_reset_reset_n),       // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (cpu_debug_reset_request_reset),      // reset_in0.reset
		.reset_in1      (~mem_resetn_in_reset_reset_n),       // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (cpu_debug_reset_request_reset),      // reset_in0.reset
		.reset_in1      (~mem_resetn_in_reset_reset_n),       // reset_in1.reset
		.clk            (mem_if_ddr3_emif_0_afi_clk_clk),     //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
