// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H)NQ6R]N95P?%?6I9VE7K2XL=:06Q"0\M2(F[#8GL>R*6=73@Q#%3,@  
HYK9S?F3CL]P?V9-+^\2V&YWZCF+4M_-C66H-5847+-IO>"Z4!W[L\@  
H;?[1B0!X\PG?R@[9GK3C(.FP5KUMB#?30E]2@#*/F=KX>_O/5S3!M@  
H0DO%3"'NQXW4JDC1WCAC^2LW,3)6RI).# ^\T#1U^?"&O<I=_7O!3   
H8C&?TJUV>;)$/D6ZA[ZN'\0].KP&O]1@[OI1>X*<Q3U _3G5?FY80@  
`pragma protect encoding=(enctype="uuencode",bytes=4464        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@W9"80UV@RP1]W;'5Q7F3]&FA+UCJBK=4B6R,>T9+H)@ 
@#;9+T!Y9E&!RU]::H-#_J^3"HX#O_])H"I)(6T> VK< 
@59YSN%S_7-@D[[86SX1,[WBQK@*D;C0)+=#=*R4+9B, 
@'"@PQ)/DKY/]_99R4PUT9 =0,8@T,DU^R4>'F3WN^J0 
@X[Q^YTG7QUT7Z*7>9:?:>RN%#9P=XHXUC$WIO&LH0A@ 
@X6LX)<EZBH=6;61'S!F3LU^+TC.C^T*]E?%1')]C!+P 
@M24!]^&N?QV?)?4W/<KA]6@A7.\%=H*0;A9^[(J^\^D 
@B"X,86Y@64G/E[+.(]:>(CJXC& &*4MC6;5'HN'-> ( 
@F=B@\:'0OGUK+S8K_&Y;&_&$2MJ:*UT1J586K"!27[H 
@,6SC19EMG*=L\%TP+@*FS!ZS;;T?MD9KE>(:J"SIO7L 
@,=C20< X>[;[=Q\7.&XUR>I/4;YGQELVNY$!F':\JP@ 
@]O3ZFN9*QJE!7Y1/N"%=8QE?2E'J0$(2B]3K,$84V*D 
@:W::N\Z]$Y#]OA-#P52<AV3W %'AH[5M9TW,DZP'DS0 
@%+76QUL)<Q9@7ITR7J"V\*TL_A=?TLWT82$QDO&LH8  
@S'X?^0<#T)+;M,%/JHY7C"=LI0R0W_T=3/HGN@;VE\D 
@$:>WL4#4C =]FUX8LXY:OY4. ^;&0O2JD%[*/QGYG7T 
@!E1X,LT9\*_@WL10;+TE#3,6NO\L'O_ (KU#5;4/L=P 
@#0))9=> -,_CT&EI7F4%_E<;I'>TNS/=F$DZ*_XZP20 
@T:8,%\1@?Y\#WS>Z&]OL:LY<41&E3=6@6.X^6"U$)1X 
@P>@I&<P3MV,(H[IE,A1BXX)?U'1>0LK$JO^\(S[3/O( 
@^<_7M;HLMF9^;A"K@$72PY7F,(IB^5W\ZF8>)QI8G04 
@3>B'8@92NL/%.W;WBD;>94H]:.3#>;O2JUBR54L>?*0 
@Y+1D\>N2<?[1I.5+^!PO%F0 %%[^BSV:,=,ZNRS\!'< 
@BLTJI\%00A##19[JQ:M&#$1GMM2UMJSS)R7H(=[IO<< 
@KU=:\0:TVXXB</(=!--4I)EWN=FA*52]$5LM!*ZMTQT 
@&$R^^O2^N+UV30B\FD8"8N)Q5R7I_OXR%P\&4=54*"@ 
@X/8S9?JY CSF5^P^*V(/:D(.[:[H*R8A2@.5 Q0"H8  
@.M^L0\@,$E$U5+;'M8DX@[KKT7#"-_\",,XUV(TEL)X 
@OB-L^ID[J&B+Q":7LPU0%78K+52HI$*>T,$([+A#(U  
@7AC[\Y=1"R?>/Q)\A:[Y)75J?.8EJ?,R7KK&8RL\Q=4 
@PD:Q!2]Z03S0H@4A>OZWZ.@'8P$M%Z<$YJ2(,%8;#OT 
@T,8UI.<)I387R=Y%.;S4)@]"]U T3=[+U4!7>\L[%!X 
@1AU_#+<_'(<;B<R>!1GD\1?T4>.*S?><\UO"Q&%-(Z  
@1\4;3A\CU?*Y6WQJV3,LILB=S \/DY['W^KR H<(K;X 
@R!%-75K*OF*&=W^FEKPS-22X)1?TYDZQ7R3CH''^07  
@+/QL$:2NZ8O4 WN[!R.E+YYY)<VAJ,G(C*8CC;C$8+( 
@H@+U)R@GER -:MA#.[#=EGK.M\G&7F/,ETZ%W[<<6]( 
@@K'VI/LD6J3".",!,&8#CFVX_*\+A&"H+#,>L^X7_G( 
@T5Y,,.1@QM$PDJ)EV8EKQ#H_-WBQ[W+!.&KT$WHX_8L 
@A;Y 29UY+.5Z"?J58[OXB+YHOH%$M/8P[;_OMNTYJ!H 
@0%EY*^D+^E 0$8SY*TXFVI*%/),&9=TI"0T$,7"%A^( 
@AZO1WRG,81Q)]K5@')X<O+B)65IYSRQ30^!OD];D+\0 
@5+DANZA75D.-/J6ENB1J]ST9UP[U.&A?>GA9M[O]CS@ 
@7G+ZVX5N^":"* ^5NR9AD-72P=(5R&X6@5SFB.Y;P0$ 
@XC9W?(+:=.(UIT?U2D]%$AV-],,ZD?D5.2/0"<FC&DH 
@IL+I9M?TDJ!QH"C1Q,U[X(!T31_^'AV[;5\B@?@U_=@ 
@;[NH^]&M8F0=^$S=O\TEE*\FC<V]B!EH:4=M,H;S '< 
@"/]8G8FF&%"MQX]36L) 834ELLL-S12"\,-]H05@=", 
@H^A\>$S05.1H-QTOT2Y0O,*M?+M\'-A8$B\:IDR/</P 
@]L$@X6.=U7<&.PCXR"FRM.,62< @.]-6J62RN<O3Z>( 
@ ZK;5?(=/WA.&= :,B?^JQ\F%?*%B?4!+4R )(5[1V$ 
@967>\4KU$?P?*T#7+_\J=HYJ0ZPVB$7;JT//9M,#2:  
@_V<T',E11'YD>R]I>T7*S8*SQE//HS; OD4%]>FYTX8 
@E_LSD@:'519S%2'DS_($P-<"NHK([:H5SCLA5@5:1PD 
@FUW='IS;UXJ0P,IZO,]UG4\U)0"X16<<H3 F.A1<<A@ 
@%.U@/:J1U-#P\_9[Q6N7:2=CP4*#@GV_,$YM8]$N=2, 
@9A(G9BT^#O4SZZ5$/8XBDQ_1'S<2Z]0CS%;ML*8]GXD 
@PT^IAO$LI*$479_B@&G0?.7GA:6MA#AX)_4(Z6E\R+  
@<0&]'CDZ36P<"Y_*#P&]?_P6W9RJ>K81$&.*]#Y?R*H 
@K@TQ^I07(>HYJ?TT'.3)-8<K@L9R43E;G#Y$+#21IM$ 
@VR.CK%C?AZ89G,JA(':APKB@&T,EZ6.IM:Y,21$O 0\ 
@27C5C Q&.S&S3,%!=\T*15SC$_0;>LU "F6P!#(A32$ 
@L0#FC;@QJL'^Z*_;KKO FU0BI1\7M<0+?*H#/>(8>#H 
@O&8<NJ\PLYA,8V@96D2OR=4R!;Q<"0_Q#+4[TATZ0%L 
@7>2WSC( .,JFD3WE^H$&/>OYX 5P)BHA8&:I6-C-760 
@61*:$?+N6DNSNS&L&5Q\,^)K7;V_O(*O@V$0*6<#_DX 
@4S\V[@^]O8*K)%"N@#EU%&U5;_,00Y(S,B(IAQBOC,\ 
@N(2P$#/V@3B1-+GW%P_N;S]:NE%#DPZC/N+0=)T1>,\ 
@,5-\S:0]=D<WU\YGXL:!0#0 397_/J&(^(.)148Q9.T 
@;6.C>08X&7)Q,$^V_<'RN+<[%=TKK$5,>^]Z.Q"P.DH 
@2Y@!OF!US0[]PUA__$G50]?[=.;W>,S3W2^D:JZLCSD 
@/$+\8B'#J.1&2<(+2L<^+NG1SNV$RQ83;P%/JX#=&V4 
@K0_Q"5<MH;OV90:YC>+GCL=;5?"&J09-1PV2I@&;H(\ 
@[?]NL-+DLCJ S)Z13QK&F0K0/14 7WC '6Y@E^%D_T( 
@7C'CM+0DFJM^+_=0<$9BT"RP"U\RCX4VS9^@)P_73U@ 
@OD(47[$#8;GW Y8!V+-V((]OCS3DO  TM9>$0-V!2AD 
@A=3TA2^A43BKHJ_D0G/N"F%S"=R-99/\Z+P=(3,N>8D 
@C5=*?;L;I<:0]-Z'B3N[OT;CSKWI((HXYM#>.R +ZM4 
@(S'F'3$1PPJ41YO<[$U$-T?&(:P9GDU=%-DETLSE<+L 
@_PD!YMTT;/+$]D8EWZ^$")?B4%([E'L(-LKBH%%#+(8 
@GA@W9PC$/6$S8E#.1R$]A(6KY3 -[Y=6P?R.3WFO[7\ 
@2@IMN\ %N$QB9*NI.#45DM?L@8J(D)C+J/_F/SR"]E, 
@4Z- OY1C38L4,)B61%+"^Q4M-LKA>Z]:Q'[#KVJ[F7\ 
@QPH4#\P]%X'-.DXA;@.DCQSK)] ,YLNZY%L*:AEC!-$ 
@YPX0ZRIHL5QR35IC\6*&1'@U_7^%'BFNWA57)1H,WP\ 
@:3UN\_>B847;JVTI@BG:V71^G)UP[:K)!%(Y(/3M6!X 
@:"592G(?0Z)"8VNCI:0> Y;::L'N+ "*4!DHN=LX/G0 
@3"()TE[E0[&.!/4M3W#P<R!T@#RP\P(:*?[7CP+R<.$ 
@\N+O6X1WB2PRN&.  ?4:V)EQ1@$0([T&2 ]Q K_UA4T 
@^ROK[T(K6$W7-99&U>&H1>*S*UHHQ_2]!0MK_TA\8A0 
@+1F'5PH,PHTGK2*;0+>)\?OS:HM4BF0/:\M0N: S"0T 
@SZA3 28>A5U&R%JHEOY'(D;A-RD)K)>L/89U4-%#XSL 
@J4335QD*13R6L#+WD#Z;IW6%]#B2[HXW4X8.)N)&DQ  
@]@S5P+OHR@"\)WW%I%AM@:TA^Z.77] ,XS%I9/DQ\G$ 
@/,*^&E[BX^_M?3<6_K[Q[&F@,YY.,L\9K"LY.RH@&2L 
@6>F][62X($@M KAV\#94V4;T[>W]Y*8H.^\48^2EIU< 
@9ULZ]&!$Y-N=N=8/7$W,J2:9)0*RVDJL0P)9O8HU=^8 
@_2L2F'.>"RJ-6:_2LH9)RC>NA&H&T=;Y:=AUTY ?3M< 
@#SK7XXJZUC*KW6$$,=6RW679PD0S1 R@FD%!5\X+>F@ 
@GUI:B5QWD&PL'N.#4$;6U]9W_/7X-GR3UV4>6JF^&)D 
@4N/&H2V)<^_5C[?Q6L:TIB]GN,W!GH*I[!)+G:.1R[T 
@$II?^+F8<337O_ +:R T9=5ZR7U6H1Z _#G6E^T(GYT 
@[0U*JFU-"I.4[^5E2W_(BP*9819*B"[YT)H1L?]5D/( 
@RLX(SK@PY20]ZWM8$]J[?,T:^F51M*F#\[)KG#]Z]UL 
@3O%1,\("09#PV<)W)S3&X'!"=:-9,9AQ:=$DW[#&>A( 
@8.I5X/(I)-"LU%VI>DH0M4-&/D[XD$=;MB0_8S4Z*OX 
@"(PN[5DC:,=HB ;DC+ FY9*3)F0*!VYOIMUVXPA.:E, 
@A.81L$3-Z0($K.@@KJE3R$;<.5'E)=TFI<-H^^?L^*T 
@OIIP)B@(DVQ@2H !X.0^?-X<+"<RR.1M+PLCM^R% 68 
@%-:Z*5,#.35Y;VJHF=" G)[@+Y?$=#TDRY/KQ.UXQZL 
@$D(D45DI@(*6JI0;*1)@HT)]ULBD F@KW6/*/>5(X24 
@R55NTN*._5EWM.;XC>!6E;K<I%]Y'2SFO6\ZG^(-\20 
@$0P4EX!&!Z_O0G$/<KR!H^4RK..:I@W$(1^5<5.TVI( 
@#&6+8,WVASQ2W[AP8^_@H76W#'OWVO#[DM)_;_X3)80 
@1FM?O;@Y>\:L9"P(K%>!S]1*SP<FI*:T@,O2U%63>H4 
@6+$ \[O4N7Q.#)21[?H7'-1L?O\.79R=LH.KW"E%B&X 
@BMWFO.68F.:L-O3VW8A[0CPGN]G FOQ:P1M!EB(+!'X 
@62D[S]83S]OV+'JVD]'\E=(WLVF(8Y1PWM/IB'*8MZ, 
@(TR/#8HE+H4GG-.]Q*^-K8I%TLTHS5\%:,]#&D[&+KD 
@Q,8O2B6>'0$:.^ O[WSHTPV?GO!,/*)!86Y.V 3VFVX 
@LA7ON/#W05,"[CLT(D$X'2U?6,]TTRGJ(*3IJ*QEA0  
@"W-_KBJ;D^R0*A:Q/JVV*.ANF;;-1*S D$Y"7NOJSN@ 
@U_;.\8KNF,8PH1R,?2/#^-C41!%GDKBQP5) ]+^A@+( 
@!B\8JJ7# SKM7L*!OZ[D/-,YW,#H-JU)>!E;C9,2#M8 
@##ZXLQE6@5:-$B2HKIPNY5!W+7Q#_?J//@>3^C\E>B0 
@@VT7)PSR=3Q#^8YC4-#\2P6.\]K"Y%>98Z#7CW#I@2  
@K4W8SZ7HAZ4\H4KT$\U3G"!E=EL2RBS?&#/7JH=MM=  
@OYP=%X#%(F%\AQ?Q6U%KY@RB]=\EY%A$][!_*SE^?8X 
@9/)M_@7.1&WB@SA;JWP>"0(?$?+LU9[#@-TJP=[(8N4 
@9>HG5HN02]^%Z4!RV;R6Q_'7U;8\"L.?V5W:]CL< 'P 
@4V!& 0J+7T]!0!<U\@/+A$XI[V28&$87)^V<J4]F-\\ 
@Y"[6D5#Y:46#_ 1JP.F446U=7&#NZ&%J*R7'Q8=,;%( 
@?L>"\B!Q#AB78>[C*8.N)C[5U_U3&P:<"-FH,68_D$( 
@YW6:J\L& ZJJE/W9Z)1IL[&VCHIH/\V.C6+'#'6L[1T 
@/7$[^:+)]^&4L*6 G6%YP+*L#N_'"P8<\?:)O\L1CJ\ 
@Z[=/+7FPKP%@1J7S#Z1YY1/N=K_>C9*1D +G*0HG3@8 
@0S<OV 8,FG)* "WOL32<9[KE!,L5I,'.,?P0ZY"T5^H 
@9Q8E;,$]A\&M/?2^C^JTHT79+9M3\KD7SXC%:!\C@UT 
@%('ADA[_LS47">M3ZZ49E#P,=-+TK#(Z6 4U)0[C188 
0??"\.Q\O0ZY0;#AY&:A&W0  
`pragma protect end_protected
