// q_sys_ext_flash_asmi_parallel_instance_name.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module q_sys_ext_flash_asmi_parallel_instance_name (
		input  wire        clkin,          //          clkin.clk
		input  wire        fast_read,      //      fast_read.fast_read
		input  wire        rden,           //           rden.rden
		input  wire [31:0] addr,           //           addr.addr
		input  wire        read_status,    //    read_status.read_status
		input  wire        write,          //          write.write
		input  wire [7:0]  datain,         //         datain.datain
		input  wire        shift_bytes,    //    shift_bytes.shift_bytes
		input  wire        sector_protect, // sector_protect.sector_protect
		input  wire        sector_erase,   //   sector_erase.sector_erase
		input  wire        wren,           //           wren.wren
		input  wire        read_rdid,      //      read_rdid.read_rdid
		input  wire        en4b_addr,      //      en4b_addr.en4b_addr
		input  wire        reset,          //          reset.reset
		input  wire        read_dummyclk,  //  read_dummyclk.read_dummyclk
		input  wire [3:0]  asmi_dataout,   //   asmi_dataout.asmi_dataout
		output wire [7:0]  dataout,        //        dataout.dataout
		output wire        busy,           //           busy.busy
		output wire        data_valid,     //     data_valid.data_valid
		output wire [7:0]  status_out,     //     status_out.status_out
		output wire        illegal_write,  //  illegal_write.illegal_write
		output wire        illegal_erase,  //  illegal_erase.illegal_erase
		output wire [7:0]  rdid_out,       //       rdid_out.rdid_out
		output wire        asmi_dclk,      //      asmi_dclk.asmi_dclk
		output wire        asmi_scein,     //     asmi_scein.asmi_scein
		output wire [3:0]  asmi_sdoin,     //     asmi_sdoin.asmi_sdoin
		output wire [3:0]  asmi_dataoe     //    asmi_dataoe.asmi_dataoe
	);

	q_sys_ext_flash_asmi_parallel_instance_name_asmi_parallel_instance_name asmi_parallel_instance_name (
		.clkin          (clkin),          //          clkin.clk
		.fast_read      (fast_read),      //      fast_read.fast_read
		.rden           (rden),           //           rden.rden
		.addr           (addr),           //           addr.addr
		.read_status    (read_status),    //    read_status.read_status
		.write          (write),          //          write.write
		.datain         (datain),         //         datain.datain
		.shift_bytes    (shift_bytes),    //    shift_bytes.shift_bytes
		.sector_protect (sector_protect), // sector_protect.sector_protect
		.sector_erase   (sector_erase),   //   sector_erase.sector_erase
		.wren           (wren),           //           wren.wren
		.read_rdid      (read_rdid),      //      read_rdid.read_rdid
		.en4b_addr      (en4b_addr),      //      en4b_addr.en4b_addr
		.reset          (reset),          //          reset.reset
		.read_dummyclk  (read_dummyclk),  //  read_dummyclk.read_dummyclk
		.asmi_dataout   (asmi_dataout),   //   asmi_dataout.asmi_dataout
		.dataout        (dataout),        //        dataout.dataout
		.busy           (busy),           //           busy.busy
		.data_valid     (data_valid),     //     data_valid.data_valid
		.status_out     (status_out),     //     status_out.status_out
		.illegal_write  (illegal_write),  //  illegal_write.illegal_write
		.illegal_erase  (illegal_erase),  //  illegal_erase.illegal_erase
		.rdid_out       (rdid_out),       //       rdid_out.rdid_out
		.asmi_dclk      (asmi_dclk),      //      asmi_dclk.asmi_dclk
		.asmi_scein     (asmi_scein),     //     asmi_scein.asmi_scein
		.asmi_sdoin     (asmi_sdoin),     //     asmi_sdoin.asmi_sdoin
		.asmi_dataoe    (asmi_dataoe)     //    asmi_dataoe.asmi_dataoe
	);

endmodule
