// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HY8++[[\<Y "SW/5U[+>CG:JV-34N0A%L&7Q15#)V'8M_0QMJ Y^2D@  
H.^@<WZ.<X *L2FO>'-53YV[N8CSHBJB3@7[V6B> 7A9^/D%6KNH9]0  
H4M<%H!?.^<5[ZF;^Z+#AH"Q2TN:YF-[J1,7<\1)1 E8%T3,;<Z(Q[@  
HXU9[Q@@(XT^X0:G9.)>\O.\--]?\[_6 G_ \4JCDUJ8.P2B.]]51@P  
H::2N\P?'V1^(Y52\H;I]\XXQ"Z_Y$N^H;PA5@&)$B]KEG\ \%!D8FP  
`pragma protect encoding=(enctype="uuencode",bytes=3728        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@CT0'W^MSXCCPGJNB#X 3_?!W,_)W(J+(B" /S9K<*R8 
@5_AZ@NFL4.=Q4,\.WW5TN"2!1A\SMC:!LT?'!)< <84 
@\7\BXN.Y0BD?1S=?F&!_8#N:$"WAF9H($*S$L.5R)7\ 
@RSS0R%I*T;\?>Y,7;<6^IV@4KJ,5^1^D'4/:K,0:V[@ 
@J?ENR?#N"3/:U F )!+'T[&)'+JK,:4FQ["55;0$\Q$ 
@&BA?2L8Q)E &UK&0!WC?_)^=$PAPH:>:.RRR6[[(KFX 
@\M4'$*9RLP\#(ARZDWB;2<L>#T.#5$_.JM#H]Z"(-+X 
@=6.N%"3-P"D;TW+PWPV&WKX%YEX_$EMG;1$EPS\ TO$ 
@BI^*E]&%A7&YWP/<PQO^M7RV#B"8U[4$*9Q8H_-JS=\ 
@VPTWU\][U/W%R8S5'\>%=1K!'(ZD9N"GE68\.+%]:FP 
@D3VDG1BP/M(1/>.!;*:-YDR<3#R9\RZB9"8G\_KB=&$ 
@H=<O2Y!P4/"OF"]-S?)#DD4;#'&^$WDU5 6F;L*?D)8 
@] AF%WEYDL1IGGQ7?3N\S39$TBX(USSU'TX?SX;OL(T 
@[FQP7EROYS\_]KO1N4MKV'XRYTG=[UM]58!ZS+(!_$0 
@&CEB80BA56(>7\.W_(_UZ!?.@ [S,NC&*:8-02Y6)PL 
@_0=!$.-+6)XP"&;"A':T70YB9.LFY23>:"H_4ZG<J!0 
@9R=S&G,GX]R0*?/#;5=I!27@Y5B5))NS%,R6%KOR C  
@=SM;1;P4-<W^(W/7/PY1030/G3>)R(?2]*S:EH0;\-, 
@P<3ENH[R*O[L%D5Y7SJ97N?^1Y1; #M*"34+$'79F@P 
@[N%!Y67.?$3A,>DQR@>VBY@CM2F#YA8@AH2#R+'Z^<P 
@&NAAXUQE/LZA""QY%[DIO%G_>EXU0XYY&]>?[0+#Y<< 
@%GS:L0[C<KA*^R*A(_R2@]94.U:]C56<49T'\5B]FE@ 
@Q>*[A,-CW&$;7[V)[+BS#(&\58X\3[43VZ_ U1O'\#0 
@*>C<2G?CO;^, WK<(C8]WB<62G'B:@OLE-L]D>-#DZX 
@839]*5MY':F.8,+D+FG&NOMG[)LA?HL@'X\2<QL/+,D 
@5WU7F"C/S5#[VKO'CK9SKS62 Q#U^GK/]TAX+)FX%NX 
@B\\BUA$\!-64R:/[]#<F1)VS%L?E\I<UZHP1Q>S!-7, 
@K5\%V^JOZL]GK!<T+5CL'^F&@E SXV0K)=V4)CW"7]X 
@ IW5TAN*3L#:%,TB/-]G/GAHN*5FPYBVP"[Z%<:":V$ 
@K#5A7\'=#FW@DZ(41!@(&BX[C,46!*XT<-;*EP.FJ+\ 
@?+@ 7E<G#'Q(O&*)KI @;#@XU".\:CKAZRMEO=QG+<@ 
@ K(<@WV"Y]@M_TL2G,6V=,?^'E'M-XX?GE0>]XOS.RX 
@\]<.:NA)0:O1%M3LT@>.U/VC4-"P1H^3V.L2UOXG0:  
@+K-W'BQ88!#RP((O!3;NEP*&!VEC/K9Z4B]&#<3L_#$ 
@5&S+- [=W_ZUS:R"%.Y["J<!O$*W]B<O,[I!P_>$LXH 
@8'/F37!<%Y7^0HONY='^#LEL#E__(UV@+&>I;9D3^FT 
@7IOJFYA/6UX(S%^TG&+&1>1V'MQZZBW)U@+K;'4\8-0 
@I!F-<D-$X.3[:[GERLIEA<J,:,.M!4%1XOYMLI:9;GL 
@S/)]B# Q\7$,9UOOU6LO44=QV1XQC.J9G2_,DG/QC,0 
@]-.<F,VD"(H H^]FOV9P'T8WM^+D0"9+V?\(X\E*T<H 
@22-\W1GICZP2%DATMJTAQ]-BRX&7C7"SA*  E@4-7 0 
@T5:P*=[Q1S)V37T2!2UA>  FZ-1;#./9.%]<9$/\0.D 
@]I2J23+I'!*GG@;L'\8!ALIBGD]-,YI6SG[$UJ>+F.$ 
@BY/Z%B%S3W&3DP$9-L4%F"6]:$+;X+<0A2\@,44(9*8 
@W-"ZYLT[[\+,X)D[L] [TQD)8@_%Y&6]%=IQ0<<V]P, 
@>-@(G4P0=5,5<3_JTUQQ .9_-4QPF*0T>O9R*0Z &AP 
@)4)37.0\A#"S_,"*)U 2(';@JIT22&.FE92U&1NB>JP 
@5!8UK%R1S+\%X[E #5A3Y'(; [J_AC00#KZ#)K2[48, 
@>]_BLZZ43<I>1R&+1F$N&DC4>J>BP"#QK\3II5&5!D8 
@A\GDZ< RIHK(7P-UFR="3B@V=#U.!#C Z+J*$9B>%]P 
@VB069M5>Z.7MH/6]+U_!K:1XM7JZ9XBOT^[\/*1@?1@ 
@$MJ4*9=3HRSJE"[I'S:+D19,9)E'_'[G9!0@?8KN:Q< 
@_/!+#$!T9W5H:=:\\\2N"A!]##J9+3I,X/ #[3#ELHP 
@<LXMD;B\/^YL10N#"D_DU-S-LV80=!)X3[\7I.MY,R@ 
@OZVT_^#+8DJ0???%OB:T$:T5RL?!;UM0\URA)?<POK\ 
@,+XI-X1Q6%-KP*! _$BFI9G5>Z/T\76(HSPIN6Y\)2( 
@5M^_<;4VZ_ ]O:Y*0]@L*:&(9N:]O_\B)<I0:(W<F?0 
@F20.H U4>X C*ACJ'O#,<$YF.G>QH>\&I.<69?9]>8@ 
@F1OF,J2(O)H7JR(U5<8J+/V>0F,_;IMRE:$OB*^QD6@ 
@\;NO[4FZ#][GGWUY9$>T( ##N?<Z@VPAI<Q.;1XRJ58 
@#\Q$HJGKW#>A-OW)Y3^IX&-(&XNZC2=6W(1ZIGHW=L4 
@W]'"?7M8<$<*4&H)(F\MJW8CY25266/F^*VFTYS \)< 
@NW/F"N9A?.$H6$153"TCL7NTP!.O0I%?:S_<DB&@C[@ 
@^A&3)Z&:ZB@Q(SI0+1=3L#L(B*/B\RO77F9 \RDBR!< 
@2A+J6.K$M&FC*9YA1.4069!.?YN./RQS0?D9>6TR6G, 
@% X72%\]&@A-$@8H+3./)C$.H\T7;J&<IW.'8<\*0=< 
@7.JB)/94Z7006#G'P&239?P/IB0#P46,+&.8I?<K&P@ 
@L>"693+.A]JDH(+F0)^'J9P+>=?U-WK:2_4(Z)K=P-\ 
@$'67S:#FYE,Z>&NR[_74,<!0JJQ0H6MN'@IAC;F#LU< 
@VLM7]+A@XJL=C=[D?@QY\DU5+L!>- 9%S5?2F4__><\ 
@*2IH+?%0Z</'$5^]H(Z8EDW3[YS:@U./]R#D7_R>@T, 
@+*^-CL^C:6-I3]:<R-?:.OSD;-NR DFQ6^KQXYRW614 
@R@O[\F=2%WN^?"K?&BL ?/V4@[MZ\@[.\3\";7L^1<\ 
@2J77-\IA\=2P]IZ[X36>&?X3!,LWC\> K%XS/9?&B!X 
@G5;WX/'S%3O4)X??EF5G\FO&8)<4EQ9BT@!,B\[Q?.< 
@FO2^C6EF4^-3V2^-W$L5=3$W6'_RFA &#ALR2H"'HDD 
@AS).QD5%GJF*YF\;FFO8XKKF;Y*.C<-Z+\Q+]R4PV4< 
@ORHC23CX7GM!8?Q$_Z,G)J($O#GKUEQ0RU0FRX<74Q0 
@9Z$NV]K21&*:"VYO-5]8 YE;*V;'/5'C2VYA&F;UBS  
@ .L>>8N"GPAK/2,I#/L;G3BK\.JV/$^TT;V:'TH9A)@ 
@"7E=XEJ(LM2G<H=A DAH&.H!RM8>((Z.ISL7WU?]'M< 
@CG(],7.5!> ].&(5@<D,4[=#JSM+D?XV)6X"8V;;XBX 
@EG?<Y,F,QR_XC438\]C&31YG0&P8^KBL-8VXC"P,&?( 
@;&;-Z-Y>64R$/.*S.3H(#UN>.EYYX9?#M0EQ:T!?RFL 
@YV15IA 3;SV'1YW#@*4)LWB>:0CJZU"-5;]_HNCS^+< 
@^[L1 ',_KX['G2@?Q!*UGI)<9Z-@BND#'\E9$O:Y!@H 
@S!DI5]Q!]Q*B;6L+<T^'P4S]CB<24NPEQ4C@.*\0_GL 
@+&[#R_>/\.J]E^ZU*++,Y&=-'@^96M_AV*#!&"&3,<H 
@1C.KN@"SI^MR6PV;Z75%7#K^ ..7; ,K^I!3JM.N!U0 
@,EM?E2R="P!+Z?(_)O]N09QXCHQS3[3,2E0>SPTZ$,@ 
@W"1QI+DM. .#O.KZJ3<"K_O%#H#/LA>NZ>7CM&ADK_0 
@B(]Y#M4645^,ZSF+$@'C4<"Q$ZH4>X$KF606OCEHMH< 
@CLD<=H%&XT=PBD6-<^J3Z3;3/OAN%'I5-Z=E#*[1-TT 
@?Z1U8P<0-BGAH0N]H'RS27L* +=.5$L5R9MT!W(@O?@ 
@;[30?E6/ #@6!F#Q;A&J>9?B)A)&2-()*FV,1?_3U2T 
@ND)+[5W+9]<D4/86%Q%A<F;_N?)Q)09QF2%L?)X4$;( 
@@=$A,L(#G+V _O@B%Q(QV>P)/P2SD7)_=5&%R 41&P$ 
@B4OT\[. N2SG67A4I;+D]W*[;F"Q,H;=4_$MET,GK#P 
@)GG@)>3%__R8+3FQ)RPY=:V"S*4;^39I+PP??HG-408 
@@.M0Q^G6PT\<F+"4]H?-:H_[L(8W$MM3_DY8O7HNZ84 
@K=!G#K=SMP:#3:A/S<*:F2KWZS%S"PJ7/I4^PIZ>13( 
@ :S"#-W=N1J,^6Q\[F;AL"G#0EA%NF-T"T8VGN(YD\T 
@U<-MZ?CXQ0 PP"MO#G&$,A1Y^W<3/%G;]8WCR>R5*^< 
@?V<;],V@_++>DJE*'MU:1U$UWJ[FSQ<7+^PJ+M4J,]< 
@ #_478,6UQM7AH-]HCZ74($_%PEETD!!^]?'DA'C ", 
@;R/]HE_Z>= H'#J^YAA,<%J.&N]F94Q$/_U5M6C08V@ 
@)B4O$&U<L\B%9*CM>#AQ2W;]#:<=T=-:]!=WE-8GLQ4 
@87G1*9&^"?:IJ$K^6PP#J6I9<(4)^C(\Q@*G$Q5RM<  
@4-&BA/K*T0TNU_SL1J75>UOM% .\/\5P)#+PR1YV4S< 
@A(VK^Q(IIA!(*C16='DU&$G #.-13Z^.B",CB;=;"GP 
@GE0AS,Y,")>3BM^GR:$N=[I%B?H8-GX6 $<EC9H>.T0 
@B<PTO0<?8IRSPI>)F,YM;OTD*6*%@B#6P0$.JV(3UW$ 
@"QX&P8\1;\^.R/T,106D8V3"68X3[%PL>!B)/Z+!5#@ 
@!?J/5^:QMK*3 !W6VD<K :=]\'$K.F!EJCE-U*<Z:]\ 
@)SZIYBJDW#&NA]""38RFK62FQ8YB(SD,8<F(_J.U%FL 
@@GU@$KN:8=*H]NA*NP?$+U.0(6O/,@IUVUL>J]3O#CX 
0O_[,$CRC'D<H#V:8<]B^Y@  
`pragma protect end_protected
