// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H/?;6H?'TY"%3MS=_UU/1E=CQUT">B\Y2V!2:HN.LQ^5PXB$J)Y2.^@  
HHX(;[5ZE5V>%/0BL2N@-.X1%Q4K<RB*-":W].W\O[0.[FJS;._>^.P  
HO5(X4FF2WAD9;R\*1UPWFJ2\\M/K*_]?X@K#8L@-[G-Z, H&H,5AN   
H4M_ SHCLH4H#G-X\(D]FIT=?C;DMI74'IKKQJV-/VI@SXPR<'H2>3   
HO2RL4/,]< U;D@Y,/W9P^I^.GT&^497T9(A;5?C2+ZH^.JF*:.YGP@  
`pragma protect encoding=(enctype="uuencode",bytes=4896        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@N, Y$ZK"C36#1S@]#='7S6+-VHM_BG=8UB8V+SBF<U< 
@_K:6@W-?(RW=AD[0,YMSX5OF#TGN5'>T7]&(M1^2A9  
@B)L-=^^RK=EQKPJ#S5IW(>42?@,%Y!"Z3H4IHY\+Y/4 
@!H^>FT^4M[SS\1-6W%XNY[4R3.%3ESL K?%R&%4QH@< 
@=[195(J6<2B'9:]\74E97-J*?LFQI:JMTZBS72Q 0WX 
@ 0CPTQG)5O<NP)98$OUU5 ?#/4FG="^7A(+IO667C'$ 
@R'01?7\):G#C:]W2[R_WI.&33KWIQ*ZH']KX="7DEDP 
@%4HPD\N=,YI0?"5/2+>[-H-0$AHRJIU_OXXDVX>W@W0 
@J^;,2!EC2\04&.?TM+5R%<&]4I?($''Z;\(/H;4*(Z0 
@5ND/%&9%(]ACM$^0BOAVBK]^\J-?K_:IW"I;Y@E0&?0 
@B-QF1BN9IG;0N.$\E?"P58N_=")3UIU#LH=7H0MMIBD 
@^ZW(OHSSU\!GG62@3'@%O^T&.9K</K26]@^;MND):6, 
@E6JV<X"N. Z*=0F0->+AAK/"-IN.DP.K%Z'YRQ/,RW< 
@ABHQ8JUT-*5.RP)I6/Z.02M$\Z;GR*B?I;XXL!:$'[, 
@ X11Y&\0=.<U!?U4!V"0]G";,'>+\@_J'I>0$-QZ[)8 
@,[>,@RKD81QW\NPER!@VO:#^@5G3_/><,GNYTR<[SBX 
@8I:K8OU#Y$3-:921 CS0KL8%E\O&>>X;(/O$B^Z7//$ 
@.\DNKFFFZU=$(VQK\>U_DBXCR*Q8#L,_QK#$;.;UD:$ 
@H20.JS0@["8;4>M/@1X1 :NDFC',DDO1ZR,$MP0XR0@ 
@\*>ZSAD\%66$ =?A%'S\%FQ-HQ^EII/:(H:5<]R%&3D 
@$]!V1^- \]:H"+$C0W.AR!DH;DYO1R7JO,3R;!)GF.T 
@ /T%>W89*4IGW+/0\D1-Z>Q]IX$"\SLNA!YO=F1[F<\ 
@L%[DF?[16:-!F>D,S _B4%'#^X9V,GGUGZDV!-J*'!$ 
@8KD.+RSB-E@,2T\A0@'-,A];COP]>WFE7=D+R[$>;$8 
@*S!WQ?S)L&2CS)YB1188@\>%<4=)5EYPDED6C'RYAQ4 
@44WO4R!S,-:O@ -[>T=\#U#GDB7,'>L";4J'9G6WXMT 
@Y-(VI8/:*[4,_YH%YC&&83#3W2SNNU8\6ICY53FX@_  
@F@MZ$P/C\E*"MZ\&F>-)\74UY&!R130N'0E)0K.-^6\ 
@RD R:-OW]%+3^=L.KET: J0BG*)+/_ ' ^):'^MRKU$ 
@;[:@_UG=CZ>$[_A/4VB_ RH==66V(D<DUU&IAIBERLD 
@O1/@I]I-,N'M*9<HJ9<!W\!YE%,G$"Q8H8'4CD66O]$ 
@NZJ1K=H-894!79PGR#;;9&UGA!\9P>?J:/I"AL$5;]( 
@BR:1] 'LW ZF+&#^3KUC@3;H:4W;$X,K0<6";%AOMH< 
@/RSUC9E7N[:DAC:JY(,5 ZRX;?,-K_^4,Q<<C%@0#B@ 
@8*=<53NJH RDX#ZN\0R\\[^U3$=R%+U<  2+8*&64JD 
@IUHZ,_D$!]IWCU)NE?#=KZE-IWE1QM%YU8U'?<6T12, 
@9EPF05I>ULG;J_5K0!&FG#KJJBFIUYSE/6)N.?E=[PH 
@= <^[R#5&KB".?35;<&?CGIV(&_D./X-HF%L-8]P^,\ 
@(?RV0H'=,P-7UXE5.:9D<&=*,$LX6B1Y<4H;K+..G:< 
@4HS:E_N4][>)"#WS>?)0DW)>O5_L2CYKG@&7@]WD$3\ 
@("O^K*$%TE'@VON?>ZPGA3'D+M?]^9,(JT%!,R)2!*\ 
@ZQ3D%RX43]25G-64^5G.[7KQIB+ AC^(PT<;NWOV'64 
@R$:#PP7CW<=#)1$9SH0%)9*YB@4E#8\YDA9W$W/RD2H 
@?F7V6,GZIH3<BVM7NZJ[1JV*[=:@_)&29XP%Z2J=4&D 
@,^(>&4OB)V#W:1>A3X'T%G$5H&'PV7\#AJ/F(LLF2DP 
@XI8&P$83T2U--S2?5^#3HM8U&I\5<XD@T]&O8>#8T+\ 
@6S[A:&Z8-AD@USC>EHA!^F+_<2D;8NKCKV*0GL2$_4< 
@Z,[BEZE#^^OUUUT(7)<[* PI,,__8] I(WQGE_! _=L 
@E>BQ?:1U?\E?ZYW#NMU/7(2R)U(\7SJ9<(MEZ,,PYT< 
@MSQS3];K1#[#*M)K[/ "]T1Y__5=WBA=;X0'U!O"QB, 
@(ZX'+_DQM#(A][<EH8GGE)\TT.:#=AHZY!VHJSX'! T 
@JS'2 (9;#J3K--KK'27<<O,'/W^ ABV/(.F-LH(-H]H 
@\  ,=;6^*YP_-\0/_^=ZK6,2L>NPI$C+"_F(C*YM<R@ 
@*&M#DA+^VM "/CX>WG&1\P:-=UV#;:10MZG079)TD*X 
@0%MBF6]1T7OC=TW074(7!W!R(U#Y'#UMWSP3?%< 9 H 
@&39L589_%R,3,609WA.J'A#53[/8,S$*K +R0//,U.P 
@FJ-HB_C1Z?86N[X<G/K]FD"1+3+QC^V_>KG\1A3=%Z0 
@I<91]__;V0C/?O9CMO\N].^ASE-;\!620 4D+)+6K7  
@P85@E\'\FQ/0\DFHE'+B$=4H;+NJ XQ"KZ?/UI4'2G< 
@\$VOB,F*W#MI_RA<D"92QC+=0?U"$%8%\%@!RZ&Q5!, 
@U"GA6=/GDB8,NCOPO/Y=:%(- 3UG*  WL7/AR)]P<.0 
@\I P1Z7&3%S') 5^DC!/6L!BI$D2\;^9K9A1Q76<E1\ 
@:M0&):VD8GP"?7;VX6K*KC37@I^($ ZRF-TTH^:.@_P 
@X-5G0U(FT9HJ9GS+EH?9(F/5LE%K((I%860C_?J3(   
@M2O^XN];1)BL_4R#(DPV],#T=''9MC$N?_V5X]%*W'\ 
@V<HJRN!AOI@X4C&U"7<+0)=;HWRS8V$#A"S+^.X?2/( 
@5$LM2(]]([B,"7#;7A4RY)L;SS;$VO@'_OZ "Y!+L'8 
@;$$1*T7!%%LQ7=2,$&8^K27VNG2%9Y?U0P\H[KA>[>4 
@=FPH*U%8$_F<)LO/YD9-7J,5BQ-X!ONR\P[/L]:JY60 
@+#ED3);NY4X2'^P.4!C>G*F28N87E TA\Q,V.MP?EQ  
@H@4=YUY5IY2-NB,2"7?+[F2*=/3P'+_#9LOCJ*@MT"4 
@=+X=M$OY0LV&U5Q_FL[KPN?SSY-\5\[9RMF5O5H2:!0 
@,!PAEQ#$M<5BH6UCR_>5'2WWX-:(=.#YISTT+DLS=,, 
@4@O.ZOV=@5:3O7:G^\'IE@I&^DES!Y]L_^1@#9BIS.4 
@\]2##:@%]S$CJ\_1,T)=\_&.1QIMU#5#.B^JL_7M-7P 
@V[#BP^M<'G!G<\@JDF;'-0LX,81I3_=#0&9!LCNZ"E8 
@)_JT%DS_N'3IL9;J$V'L\8=5XR2O=IA?_#0W5YN/GC4 
@9SGL40(BP[(;*'V9 M"JU778$[' >I5QBV1=K.X"0?4 
@'V//_=MLNMX6*V,F 1)$5[8BMDR;TGMT^5Q;,T+WYO  
@+$A<UM-MZ .GDI;,9T\)H[[$.^<LVE?1U?T%SZ+U3=\ 
@JJB,REU=6@*),3_,=NK["RGT.<#6I.IN:4Q#J3E5TF0 
@\_S4:1=,  ;!7]&HLPW<W=OR5]ZZ#"0^0J&W+0:Y$,< 
@%_<4[/P0+!_AD/U\QG7GX%!40\XR;RE=SX9P'5GG3V  
@B]$>Z$.](/F-TQ'32?Z=VP(I(6>Z/ _[OX/>U<#W(6< 
@//2D,@6",D0[.L*_>!0_M-KVHQFS[,Z1A='&FJ+\Z(0 
@L0 /A5"8%Q;:;E%.-C-&:GH KBB Y&$H.7NONC@ ;I  
@H-_11<>F&+9>: O3=G:I.FB?Y3"#^V]I$$=T/83H$', 
@-[YN%C,0]6P"N_D-M=4/V4+-E<SY"_K7=0L%MQ'5_K, 
@\ 0^'^>D!<&>?V,E6S>]V]F1WJ.Z/B@BGN7,9/[C#L, 
@\'"!3S"7UUQ+HQ<B1]H1_1;<28JKO23L2Q&E$QTK'2T 
@_,\2A>_J"60LIPIQ",0!DM U$80/2]"@-GKE4M)?C8, 
@[0UT7I-\3R)(6;*[8(I890DKG3"UD3]M/::E$UI.6?X 
@-6_)?91/W)$.1D0(KAWQ>54 SG)I%XU&PXVPK99=I6P 
@0^;N2;C\EF5TDJ6NM1_3+P3:K"3+31Y+JOKIP:P<FCD 
@2UECNQ,I\1V5:<9YQ7:8(U+D>HUL+U!T0BVI7B#ZVW@ 
@ [,/3IKYO%.KJ'Q,=8,KNDPR4X%'B10](RF(%( V) $ 
@,UN]*K7<F\'6>-P.$-P".B *A"$X+CPR=%'1NU/?[@( 
@PR@_[>X:%20T^_#CJ<&#")G9"&* L7=8*"D[G],"9&0 
@!,#ZV60+-7/L1M'-<$XE3<^61WS@&0V17P&#9[<*'MT 
@+$<KA/WB[Y3%\7+L4*I),WLB(4P;O)/BHUW(WY_4:<  
@2H Y1(I65UV5B?L5^*',ZA*+1+&KVY.=WT@+U[Q/-*P 
@9_"/%@9@3O.?82=#*$6Q\L8E?5@MW7",Y!VKRW4?Y<P 
@ITXA!;(VUX^/"9QO:Q5R:K];!%\?[D[?Y#=!K-:TA+, 
@]M]>U!Z*ECK+?A9BG^=UP-@^>+@RZ]V>,\T4M$&6>?\ 
@V_>L84'6L&%L1DH[%29M;,T><ZN:GX5D3<VB!>SCD"0 
@Z0+@D<;BD8]@PTA4[B[ZZ-7-V VG$/5'$L;9B)RT:P@ 
@V!#Z^\\23&L-6C<"#X]W,S=4Y3;@N+_+I[9\1@'+Y@( 
@]:,%M6S# %#K6Y?;]\'IW8SF+%:.Z<76;O,J4CL=N;< 
@B^+RA-;D40:H:NN?T.8F!30171HORIAEL,)ND5NEW4$ 
@X2@;K10'?/28?1,+:\&Y:$SC3^55\R7TCU=^*<+=Q<( 
@VKY$V!#WF!XLB"LC+OC.!OCQ-G: &?M%:K_*8<^Q8OH 
@HMA">B-PR0,F(10S0EK,';UF)SP[.L]K3G]F "4Z#AD 
@3M$W^[Z/M2^01S=FN,5H8^,1:/T53I,JM,(@Q]2F8QL 
@X\;45+@$INXN9W@UTO(HTS;D:WA"&32G[_OB\[?GXY< 
@$3?UE;K0H1O_DWB2A10O"!U<%*\F+WV9Q)(LXR"%QN, 
@I4EJ%_/%-?_I#:J-.W:F<G(=)Q@A_IE)C)-X$"BPR.$ 
@T=K#OX]#5@:1A=/DP3W]T+J@SK%&!3*^R@U.C0WZZ$X 
@@"S<C'8G7U&P,G$I> "\J8(+R<J\%U1X/Q:%X0@#,7L 
@,DKW4HN&Y_QO22"A8!214-5)&-IHUUT)90D8!7=#>F$ 
@2+R=HUS0J9.]ME_AQ["J/CGNOO0B3!I5X<#5NY^UALL 
@DY_>U$,2EOAB>+A$7R.%$BTYK-3C_G*X=G <T4@Y2[X 
@ /G9P)H""S-0H:6K04GOI)%Q=BB$N-K/FO9647ODP10 
@,/2*O^;+4<+]'J53J)>6JLS=Y)G;_C+<ULX;VC-J;(( 
@-%Z$NE%#0O@LZ66R@/R3D1'&0A"NX%>LDETDWD8-&^T 
@P_2SZ+$.3OK4(F/=E<<]2#A) $0/UK-]'_691YF:QHT 
@KT'+;/RHDT&Y/Z!W7[HF9.X*1E??T'.#R!.*<EDMB=X 
@$(N(N:!V:H"S'>^WXK0\'IMV<F\M8_!,@,:SV$FZ[&, 
@V 8#OWW#]X_Z 6;POI+3$_L#*MCM?L]TMK?;Y'3J\48 
@G]]#L_/&"0\LP$+4:R8*_AET+QO@YW';GQE$&U3\3?, 
@B;<#"WQ,N\:JFG0?-O&/9/<OSITTQ1</8A+AL@C>;_4 
@3 E ;(=_M&":HQQ;2T'B4!X=^ZW6#N8"ASG*6_?T4O0 
@7X*IRALG J*_.UK P':8.X@5A?P%5'M;ANCZ>:>F'D  
@?H&7U1P*MLGOI.<IL^)B>'#BP$+_30+ 4U910,X9R+\ 
@4<1@K3_-:DC$*2:'IN$(6]#G7CUHO84:*5%\ >Z]'OH 
@ 8NL]!]8I&H4EA=>H[VF%>?,B@!6Z:6>_ONJ:3CD 80 
@NB@P;&07.?]:#Y_:A5F@*8F[+9&R(IVSW949WTYX2Z, 
@9,4FT@)9*T+FN^P03/R@[RF!1>U<_-B:9; BYGDX6N4 
@ROR2'(+%"(TLUQ'W>%I*LZF8MG%+*/]U?7NQJHX,9*< 
@I^55?O2:2BB@&CGN=(%PP*&I_I@$+PEO'Q-M!4F:2H0 
@P*Z;9:,:_,5 *#8FYH90H>(N_I"3K17#^<J.40XYSQ4 
@;_E %2K2F; ^ B['OEQK-$K#])(D>JJ61WHWFX58BZ8 
@+V5&(Y@;-FZ\L2PO7VY=#.UQE_ SQ?DP1&F]%OJ4YAP 
@YZ*7/KH."\C2=:O53H6'_XO=/CA>TZ3>T#^8HB>HW_( 
@0PI"NAIW?A_W"WJR-)4_=BX6BO7*U*$CZ7S8AUNH+[D 
@^EU?!1&.0V:-'F9L52^0Q5Z;NQTCL+X"IO:1= L4G7\ 
@41M0@M"D@8W*?*<3H /%@9J3PVTQT^JINJ<'I>C(R18 
@?JZ'M^#2-+M$0MU@I[#!KSP>.V0]_)%$8&G:."'((G, 
@) .(2 -^?JL;61Q3))"R>LB*F<P^,('KU=%XJ2*.P", 
@.'0K6;PEM6WFJ6E/-3US:#;V^>4$KA1>BMU/%N<>>9, 
@P-)BQI)1'F:<J'84/8+-'AMRXL]1G>QU'A/SWI^R M< 
@"$SVK3'-$42(ZG'XOLK"(,';T1V=M]J6PN//DHS;0R$ 
@,4*DD5=87S0!&#$3$4PA.+O+3_?:."A )D&-09X4+KH 
0*HK[6.!R[(#>#\X%:&ZRH0  
0 G%*)$WNG&ECE;N&D/@$&P  
`pragma protect end_protected
