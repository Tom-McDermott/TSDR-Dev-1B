��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�w�����)���F�+�L�=)���ij(�P�q�����̉m�{�E�L��#�(�j޵89e�Is�E�����ߨ��A��\��ݽ<IuwD�Z�V�,��_g�C)r谚gCc ��#�����JM�LU��[}���Q��p$�!�%������Bfk��t5��4�S	�頲vwK	 )I��sL��tv#��:�]`�����$���r`����YzZ���$s��5��� �k�@�x�K+	%��p��.?f���2��}
-�<ߜ�Y�~�u~D���Ҳ�&/��C��W���Λ6�뜃[F����O;���0��ˇ����xs��C��C%_7��6(�l����t�TTk�Ş�L\�;�Ů=�|�O,�9�9ۜ��B�L`��O��v�k.�c�D�.S�1�me/])���`V[`�<l�(.�����>����s�@��۸A��W�D��XY}Ix�=�{Ry�����Z�`�e���9�W�L�Y�jd�VjT8Wg:�
�C�d�#��YL�<�r��2i��7�'TQ:84�c�f������P,�94�
4 �ꃙ��nh�GɀXMNH
5���A'ň�z��?�c�>�du$-��O�;	�\];���B��#����l��r~��&������C�d3o��)Z5ǔ�zm]��N����{8�c����<��P�u$B�!	,i�q���	�ޢ�07�he$�Cm7�>���_&X���c�V���%o��{LB���M^��1���adӈ����Gr���*�Jd�R�gs��o��74}�t�+��n��������z��մ_XsP���4l"���U�p��4)���e���&��~��C��+~$H����;��e�Q��c�w����=Y�#��.nz�P�5�j|tn��kQa�X�}l9�`e{Df�ڕN�b#�y}))�,Zک���1�Qt�w�Q���Un�i`�����a� ��7�w�_u]ܼ3D<�8��̭������[�΍�.-Y|��(�`"�#B���b䅨��Xp2�c�f�)����)Ct��$��,���f�y��6����؁�W)��Λr'rn5J����Q�\c�E��O��Wd<"k⹱>��SIUZ��/�����7�*�+�0�=*݊�Ɔ�l��_���]�A6�-౟�v��V/F�.ԴѫF�v��s�i$�+�/*���Z)���Ĉ��w��p(~a�璀Y�,1ab)�I�C�p:� G@����Q�&�^�"�,�Ut���"DF���O������8a���Ȥ�)�C�o�?���c`�`�.Jp&��ۑC�$�e�������Vݼ�Gs(��h+¿ϛ/��������*���9���{�s��%IǴNqRpXf�����O]|��p��h�4�W,uH0�A{+���� ��`J>2F������H
4� �7��W���*{�'_`�5/GT�A��Wޣ�FX�F�<Um�:)����#��&L�U�K�/ԊJ��$����Mk[ ^���٪�H���nZ��9g�N�M�ki�P��x��Q�7Ol|���s"��� ���w�|��c[��sg�[g�f�,2�A�Bj�u����֘��{�t[bW�MS|!��m�r�����B��w��������~ߣ	S!Da���@3�X���t{�ɖ,��d�tc�U�[��TOD�������:��*W��/Vv�k/��u���uZ�ӹ�AJ) �!r��h�!-����%0�g�셷�/mzB']��m7����~u��5M�eo�h#����2Sc,n/��PBD\������J}�5��~��E�|�a*z�:�T����s^/�.fIlpX�?�f;Ցq���~�#׀��-�!���k��Һ�d_��:�"o~��1���l�dOe�πa�ӳ>�C0���:�?#�of��U3���b�`Z�;-M+O
��~u�����Q���h�B���Jh��ۃ�Y�}�4���>��K�>Q�Hp��C{6>hB~_�>:����Yd��*�;#��d*m6�y���r.�'�v��1gp�Le��:C�cc���Π8K ���9�9�Ict�����rFu�^:���~[�S0��L�������f�W�����MطF�����r���;&�/̇�1��,�Ef}i��4�6�\��`n!��Ȩb�wi�q'\ ���`eW�4^��&�"8�������,�H��ia�N.~#�����)����m�zH@�d��,Fd�2\D��%a���FC�?3��ov�W���b#���#B�RE*�GcA�"�a��8~!沢XZ.�?�mv$����W�d�;�m��XD�ߦ�zϽ��n��zc}&U�{�J?�\����->�Á�bÃ�L����@�U"�^&���΁A�*�/��� c�b�L����n�)!�������г�$�#��X��x��V�8%��;r��:�z�Ԅ��ٗ5�ǔ5�4y�.�Bh��M,�RZ�jD�7z궳V����[<�-�h�fK����/���1L�x>o�Dz7O�������H���F	;;`���U�2��[So/<������דY$lĸ�\,3�E�g��O��
��ٱa5�QY0� J,��_�M���,�*&,'���o_)�GR�;B��!u����ح�>����Ӗe}�/����*:.Gf޺k9�����q�!�6ꯏ�[�1C[��y�@	l�-���i�-0O�^Q~��c��{̼e"W��&?���� �~s���ѣӓ�ʉ�h��a|�4XA1����5�cD�8%�׏�_7l�]ύ�aJ�8#��?�x�@9�h��A��5�nL����	~�������fscn�kZ������q�!�<���@����u��G�a�oeO>ul�tE��������v&W���tZl�	hܹk�'��w�S��[���r:lR��|�<��b%��Jh��{�4$4y����7�&H��~��&'���Q�ZK�sSm"ˏ��Jjњ���Y��ښ�=�I� i-J�@��ه�;�����@d��_�n�$L��dI��:Dq:QyT����oq�Լ����S�}��/a�z&b��; ܈��zçctI/��U�)����Ap�=}R6��"~ڂ���g��1�ÇC-����`�˚F<M�V̀"^n�Ɣ�h�c�o�0�-�Q�M���5��.*�Ni?�>ǧ�yS�T!yS�UN��L�Y��Peh+�y�I"PR��1�vD$�W�G�y~#%�Qu�'^��3U�e�'�9�q� d�d���#�0&��n������jE�	ǔ���Ъ�ܖ����R���V�/g�':�c7�X�s���)1��P���
��1T, DsH�s��.�GoD�#�apCg�����q���jX�/�h3�Pj�`�h�~]n��d ����(UE����r]u!�*Wf�2-�����#E4�������OkDd���Dm��c�C��w|E��:� JSS Q*��P���S�/À"h�7A]C�Z��̮S^�C_*=�اg9�V�`щ�j�����N�]|Rz�ꌠ���)�H�1Sx,�t<!|�����Cl��/����7��W�&2Gh�-���8�>E������/�� ?���D�.IVR�O���|�, ��<��8�e�u$�����^+}3,}�ȈA��_}�c/�Ҍ�:M伍�	� ���e	"B;4�������d��9��<���t�q�y�!a-�&-%*}��
9bG����	�#����-�MW5��-���]�%0��Ӄ�f7d�U	
���`�ԡ�Q�4V�{����ĩ�6�gِ�[yjn��~0���r�A�." 8�ӭ_I#��}K����f�MF##���7܂7_� �<w�ؚ �Ÿ¢�*�ܮ���Nwij�9���*��X�N,��Mu՚H���T����M	|�������3Z�t�����yu���Kxl`����89$@���}�=��ڜu�b���Ki�5�9��<���YA��x4<GX_;�QƳgE��qՏt���s�o�kP(>v,�-S���Mnf��!E�~��Q�ϑ��N�n�U�rV��m$���N�PAfx� �5��p"+�">�����B:ŝ�p��k����&�����t8����L%uPt��R�V��J3����<���O$��ad1FH
7��b����˿��C/ ��	�=�^$	w�4eL'c>�!M4�Ʊ����˟��O6ߠ,^�Oy���s�ba���[	^����sP�P��I�;��gfK5ɦ| �$Â�{����!~!.�-���~��c�I;�ۂ��<� �x����06��[�7,:����A�n"��X9��-d7��C��X	��gZ^WZ|�4&�٣9�*@������O��,��ͥq֕L����y�v~��9}�DZLl��<D\	7�:�iQҡ������$W��%�w��N�"���G�WD�!��!�F��ڞ����!y�E��m±��}�3=�����o�eӈF�P�J���{& /�NG���ɠΧ��(`]��>=YpSa������v��Zf+^uw-�d�^��#��RLA=�4��χ�����AIz�<"��+ε^f�&wzQ!��K����<w;�=)[y�>�K1��5Z��8=��_Y�>��t��jC��\�jC��
09�� �d��ğv���+�ʽĜ4�uR4{�S
�Ɛh�3~岝�ǲ�ɠTv<b�����]�1�߇t�˻�p��Ng�+ੀ�6
�9̌�Q,�l-�MMd!a�K��ͩ^��~.i��.�L���k�O	�V)� ��G��dt	H��x�J��5� �\;�J$%�+lI�o��-j�[|;�T ?�\�@�齊��>���|�B� � }���G�F�� �;z¸4��C�Hh�2�3�Hʓ�9�F�'�s��4�!֨�xנ�@q�I�	��_}<�`�ϸ�,\�f�F#��5Ym�*�
�Q"�P�`��A�����D�L�=���ʠl�;y���o�Ge�����#l���%�of��"蟓�/.��~{i!P�^��vR_���������(_�u�+�
����D�/g{E0*cl�}�G#��~�X��S,�2�g�bBr��Kv�`��)=E���ާ��0q��ϸ���9OH�zZ��U^,�5���Q���Q����[��3b#�<zD�t��j��9m����C�W�+t����0[Z��6_ZA9j������iD����MQa\� ������ߝ`�bJkx$�{I�մ:�c�p~J��Gf��q�ݭ�CI�Q��ءܘ�6���-ߐ���0���(_��M�;���0�ˀ����3���z)�C���;�ݟf����ˇF֟h�D�i6Fb�ّ)�}�8IL�Bz��񣧚ڰ�HQ��S�`2���B�P�����N��Y����c^��	އ�MO�