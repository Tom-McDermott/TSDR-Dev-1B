// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
AHcVkmQAutA+LCiRiPXRpJnobPzYpDx9StaCC0VAcX5CWyaMQLst7BiizlxG5GuS
DcJNjrca2/qa0dS1oJx5JXNFaN4GOyDvGXjvIwge7A9k6LJ5OHNriRl/BSBmUg4c
82PGg/wYe1jDAnjFN1wX+q5IbQZ+GcdmtxWQsGjEdj02GrNeSXdifQ==
//pragma protect end_key_block
//pragma protect digest_block
aeu0sTlt6akvDezi37eZnOTix44=
//pragma protect end_digest_block
//pragma protect data_block
eblOd80B6fWSOjPh1ARfN9/g8fhFmHUS++SFQu0LtZ+42l+UpKtcNureOV/o0BlU
v6DsSn2xrw1ufE3I13OXP+KbfyNdpyFv+p1koPWsGO92HwrHbB4osoFdMKECaOjL
hdFHHPoFFjlsSU8wmnguL74wp18qx1rRLZLe0xm+cNRbR7/RAZg+WLi+9FEHk3Pu
JP0z2+MyP8w9IR4Oxie/DINkga9osXM2uIEjKL5ZqdsT12rFitDCnQGH/ojgQy7A
J7VXa80QOMygcbR+eToXWZfog/OT8VvnXPuWG25eJu5AzjBAoli8qJecXiYyreFs
CPTbyXu3LVbmnDrTuhYUhmvnw7Tfu8ZW+OekhAi+DSiWc4MwpcLLni3wfEwbJgxE
69G5tiazDxf5LErRYmI/UOn3h8Is/y7hHraFWk1EAMpXEAz0jvgmb5JQm1SOXg6I
7ezDzxnBrryigFIyhN7/RSteN1W40aUErWNfECxsIS5ZeoZLqH7+ojTvUofCA7dX
vpndcDYcgsJe4Jdlg/1ANUZ/trEiMaRyYTcsFc4oSAOm4NxKGXHpjL+PxE1oFIWa
9clSJiobPMv1xm64JzQOI9SsjOVLXml7kLdSoXiz01rqprJt18yz4n3gIgIqgGov
pyb58geOBV+LVE8I8oDssZJT8MDMD1GGD+VZoZFAPqMNuc5chHOEKhX3Oi35P9AN
QiWkyDbfMxpMtQVmW+T0T9jNAbVIayeDH2r3OcfFthwvaPhHhNTAU9ogLVJnmpqN
1Y6NzP1MVLFaOSmbxDZjVHSOdwRKJ3QDgLlRChywiAWWRGhDsIgp/vbJPNWrKQt0
A4F1jP6zym5kMX9s8jULkpcfeY1GlrwQblcP7tuBY7O0br7PmO34ZZA/b+r32Wg7
ImTCi16LwfMW4IMLHRKT/92shhwI5CNKJhswEM80pxM6k8gL5qdgiBDVmAtoMNaq
62SVvkgA87ZXkYHeEM/bb3HILvjjWluD9LMtL20EfDj86LiLtQNP+TBB1o1S+FLN
MzepSToYfs9Hn1iR4qaiBmEB9/0f3l3NXoXoTUkgyvXMqhIGVlfE/KqKYhGCupIt
N+zoHYOWFOPgLqgWawK8n4n+1k1whF+nCeenSOVT0H5yYND4qbmEC0KDo8l6MfkH
e8ONtADI1FW6IiKpG6/dLG27eXKSv3LIWhtg0QXyB1irqQAEBlJpJCL4l71DyfKh
oku+6w4ar20IMLfIvXPHVAT7bI2BZzhvtNkwIn7MKqcSTs5Kof+T+4DoY/aPcwtL
7LVbpEYW65S2N0X0QY/HeSm/Bez3N0Z20jj7vwN4rWXnVNl1/OGU0b32/cBcRO5C
MZUjLM+56NTGNBbkB5eDZyb71rE0vXxpWGgCXBsx8s5xdB4G1ILgreg9ypr/BldP
H92NN8lMnKWVCL31PevvXQt/58yAc0CQc968P7YUk4cW3OUY/blvHjqxLBAoFGZG
J1JiZleCUiyHi1WHqEh5ymjwv84MhTNFiwiM0Uh1Zf3IxqyMDrCCfHYY2ey6qwUW
r/8coAagx3sftr6QHqn10B7symROaSur092yWYIi5Z1+vBuCEHhesqapkrDrRkQ6
u8KU1UZi6hJvNlPQqjOT0WJNBLfxuxcOwg7+o2wUmPMwMNko5X3ov5f37O9cE6If
mILJ1S45Jh4Bk1TiiL0YyOBNARX2oHSbV6AdC8AOg+6gGGjBk2pL20DVrkM1o8mh
5cLgmpk2RRWc+HlnZMw3KNMpX+TF3KM1ivAVkjt0c92qO5HJsq5X7xJ/D7tUBfgm
aBJ7pEaRTgLRjQLQicH/IgeJmC91BsNjfYOHUL4+rmOPH74bdr3JLqSnh9qPzCdj
JlUUetybUyah/ipS+fYO9vVrIiCg2hfVloVwiHWZ1Sqfro5UDGiS3OKqTftTE2hZ
+I4efN07HAXNfcUOXADHqRYGYzBh+UtwcH17Jzz7W5lLTEVQVEYzUaqIeujU3Fof
6Tmdy4NW4xwTw/34oqZCpGzUzOVnIQ1bYKEFBzPfPFzSDiXez+nkP6gZLMlxEbbZ
hvjL+/Fyz7v8o/Lj5KAkwCXVKrO2v+RFK17b7bSBj3+7lF7GgUo9c16ILqRmvPYx
VO5SG7plHH9BCIaq59k/+4S/LdE+BsRmbu066TLq1Sq8xt5LZ2XdXFPvelJgKxqy
JoUQL9I+dOxt/esSva1S2slRNgAjq3Af+elRqLX9HKKsnl81RbQc5QJHQy9uML/d
50r7tj91SDaHw5b/OCY2HwHPKHtrJXBhFehPU0SzipciZWfSOyAukBu4ik72vANH
xlojOSxOpeeDekpUVNhjpX8VyRZ0mxg/up98d1E42PxvSZTU1ntHyseyfgClyD9W
CV551lzzDZSBdx1mIxx4Uu/nde+dwmCYLbE5WaJbAsUifhwShWxRl9rmRMfNi9yW
rsq8Z4MJsGzUXAHZQxWrSPNtUTxD9gaKrVrJ9P294LU0mdMIt/eMv2PLiGB7jONS
mDJlwBYgRXuAj3epuS74DxSaLIE5Gif9dK5S4V2lxtGrmd4vsdmNGpr5BocolO6K
nLm4PibRanpg4Ad4J3v+MAQawE6DV/qF30SpSOr3Y8xpOS8EE9gXy4KIhwInXmjd
qBoAMwV1laFR571yLMagMg3UuWDTdQdKJ9z8VyauT/4R58eHL8v1A7UilwEkrV2m
knxlV+p1o8znuDoRba5zR3TquOiy8NGgorNtOkfHZs2NNGzgOI78mjtXA2nuuofk
ENbz8jKcHATd+BjSZJ0TYkO5gjXdTY14ABS0jv7ogVCPkPlK1KKu/eCVIYW1tj55
Jg8oehD26BfxG79T13fVGfH7A/2xi85ZQiABG3Mglp8LiR9jh0gu/ZMlpXCxwdB2
6usOa4mIc2NSP2l03dx9XgHQS0qWglo0dd/23Ypfm6jE5wC0fD+TQufPe+PNgmqj
sOW2AhG/rtHsqsYsUBM2P6ue+hPMOA1v+Lolmugco5ku5sp2vWwADWhVMfBB77zA
mwsjfsgk09EzEktdKQzwyin6p2LMSDFPd2xfHMxVpVWQhjpKjnrYmvoUumx1QKpF
E9wU26+0sxGSE3K3+NamRkVvOa2V5IaZSmZbYD6K/6iXp+wa1J9Jgv/UsGhRXAdM
ldCz5ZatPNsvMOAxTvnJRgJiMKIzRXh1dpjuxqcrOxa5AKPMrWbG0q/TuFYnLEl3
OlwJCUA2/vCESyivD/kWdJi/lLc0stDt4XfqHvJa3qw4Oiy5yXsD21PrMW6isbdT
6rAO/sLqmOqaGnEkI/9LJ0rTw0MGWWfOWMiWd9aGC4hpoID90xAu1PaDXKSWE9IN
EicQ41e9AAUOGjheE4tUTC8qKvjWzcjMJstGgy3GXS3MjIKbtcZy07ziFKHZfNlX
4pJQ3uGnxpJFFRN5dibwq3AOXZZJ57Cva/Es/yYyBjUcZ+yIsxAkL5NzCXdZ3ZZj
UCeKibCDI0MqcJkZmbFdqM+etFMTnNpWCn2u1c6HAGylEUrDK+waBLYLsRStxC0A
DEK/SHSS1xXk2fUdVcWaZpBEMoDzG5dxEfaoAExemf9DI/mmeLU0tdu002vB55YH
bBLMVnPu+m9hVA8E8sIMVCRhLl5WvP35sBOkCWCnXe3TH7RNLOG5DQU7fErFypud
d0bIFO25G3/cGK/w1T+4P34DYrujOwRPySMWQ1+W+K5AV+dzBJ+FZYuhVpNNzc/6
8990FN9iQ4IVy9bApKRSOK7IkQ3Y83KzRoXRLjFwt7YnwbvljkF/mHRaOt72nf7y
ysNr1t128yQ7N0syRIvIXJdZdjtvXC5Isjudr5Yb5R+98IPHeL05YcefjuG7LAvM
qFnrAgIpsYTdCAa0pPc9Q2zxfajbWc7c/HJU8wXBCiXNaDHXVkUnNOURfMjDJlhJ
xTPI2s27kRxkV9KkPLJyq3j5cbGhpnKWoizM6fYnKsOpMlsa3vNpCPmq1U3Tdyba
Qsef4B2BZ17bgRoHcTo3s9FWIGEUaTNwH1rBrfDgHqmpzATkOoil1Cg65fy/rCaV
MKtdTR36GmObX7+Ch6zGSAenTIvTti+8Uw3uLmbqlkJRg4nVww6QXWhRmviCKfGr
zAX2cHRP8qiJUQmG3/ZdtcS4Rd5aLid7QQfUP3WhxajULHP21NcXhhv1Hkgo9QO6
zSuSNgCnXSZ0FfqoYSH8A+gbpRFucIA2CVa/OrvBojs3MrptTcB9+f/mPYFSQD8P
v2u/qilx1o+t6RpYD13MAu4tv/rJt55FmtJdae3Llfml9fHENWRHrjdxAwh8yWjA
fxhnIFR5P35a+O8eL4BgilmZk36TwBZxqhTY7BWfFii6SWGxjsfm6spoSDLJ84zw
uCdAJlo14SM7oKT7zkHxn5q6lJNvJ5WrbR6tcFw9JzBILEdzcdK7v86Oy/S4GZHX
RacXwd+2b05w8cQ9Xv30Sunodcvol6UwspwIXDlRZgjl+ZoOJUsTGc/9bRQnblLn
jUyeFj5EzvDCwIqCNARshBm8KLD9Z3HgNlamJSH2RODPcH2hrxUcDX64kv+LaLAL
xiZ8oGHLTKw24vwjDMp9+cWm9LfjYciwBEAXPtU5hpVrpOjtQmbJzJwx7kB3QJhn
GLCEMD+92zZ1HOSOuQuIKilOoG5gXEi7u6l2OzgkKqMS0rccPImmQkOoPZQSXKeg
Z5hR+jELTBpAjPjsL9fvGc6QzykHXyc42FhCeExUeSBN2uTbFfBY6pkGv0iPUThz
jpnESs0W2sgWApUULBaJvOyn9w8rtO6Hp72vDGBAx0MJVTNuYDcqk9cYb688k3aG
CuOcptbTinfD5t5JAvHfkD1YXnzAnu0Rrx/tVSL63wXfcg5VwYA8J5qNAH8NqFuR
DKn9XW/WcRDQZuicBT6tJjG+hXvVfUYxEK3n0n3oQDuvb9f6T2BqnQ6QF5EM9EDR
D9g0hHzfBqyZjfUfZU3JNd2oEN/TIA4ts/2CU2639p1miecZgSKi32PYMKAoavXr
N9i+qvwFHLg5c1dLpg4SATZ/WIpBMWnwgid3eahZ5GvmGSIPFdUAHsm0pjRqGWus
6/zpgt4ZGeLLB2ZZjrrQaWIzFSDOF+xbYHh7nzY9YZvc/6yNAxic+tDn6wzfoung
h1n0zHrHQ4+fBioilZ1mFnFVSQj1oIP4X8qNkSiyEKtJ7yJS2hsdNtf8hLo+IjjD
7CP+7X3Fhjc+ZeDgo5lSp0tEcvHRdeE+Y4OaxK+QMSloooObPlXEs8gfea8KIzVF
nDRQyO2e4rAnlMR8UEJwBEQYKlbKj3a5HEc/W0aYwuy+foC0Vrggr7mh1SqYyIAv
k+pr+FHPvHe8yXVp68RP66rDXkQO7p3cle5P7EW9Bn9ntl9YH5cvI+nGf5IjMz/3
seJ99SlS55I+Bt3Qxsa/MKjGHPYJk4xot1Z3V1h+qvQtlaU0BYPsrW6wrSW+KQmH
pr77NsJEMmDT3T0N+BrU1eof+tb4Gf3B9bkVERRuilN53cac7ykcPPS3L0kYt/WL
jzCdqkkZCQWRRG5jtD3fF3s7D6HZxjRgpUBwdZn/XAHWYnRVv8YITsxWx7OxIUQB
ITKzrL4NPpCuuBhICW6KZZBHCJ3Nn1GDGJhF7/eN26Y1EU81YJ59+MvcmgJUNwsy
/WPsXmEVgFdyQhCR1R0D2Gl1h8Io6Tg8qCnQKiGYh/g3OXljVh7IkFIqpYJJwU9t
rZs/KUoRfHOg29vXKwy3jFWfLyOjLQGMlnplP/wUfeYHiGOyiT+k8RER6rvP6XTl
wH5ErvvczhIcyZNAxM3YH+l3UV2tyUQ9nmwL5g4Fhoo3ULo7rEPYFkgJOHA7frd9
ffmwOk4zFbCWapUuFA/JCrR8VZSPGieTWNT1i+YkNZ8PJrfXrmUYJyaC9HZHHrcp
cwwwhWzEj1+HdgaKRCIDEcxpl6EEbSMaul+OIai8t51iTN2PJmmk4QcxYM2v9hnk
Dt1ArGHgyVFXX+VJ1bi20Zau6MoKWS0I8KFgLIUKtxDZHE0goF43W6Q9X1/PrU+w
+yMEUe3BA01K4M+Z9nClEkU/eNeb5jJ03Wpf3cHSNuvuFQg8WyUZkaB8pgfmsXVS
q3ikzPuG6KpN7nG3LliG9ryWmBYG6g2R3EO4US0iGjO/UYzahIFTiXSDLeqdQA3U
zTq3gBULgdIBo0JJVAM26w7TWof/11yQodIPfp8QbQpds/X2q8Lf3FuF1YK89fvY
eTIiTLEHQernw8zz3tHlA05HS/PjVZWnwOWThzjXyaSjJAoUNFPziwYUsVCsjKr5
rvUAV85hS8XnlhAHeXQLxaXAtaTT6/iOgs0EA79pwL7XnktLfmeJURA/rJsLRSkR
5UfBDXuDLtMXhOsD0ZdGhCfmwPsEv5SEdcslRYgIt1PWAT0Ft53UetRWOOnIOhxb
LtFELHdASwsl6Z9vZc83712VygBVV96tTFgwk2cVp2VVrVbX5R3qMvWLEM4jAev2
3LSYNUQVZ13z9BDrwm+6TCm08cTYjozObX7J6EYHKz/pk6ZxogmYkUTXV3HC4UqR
5/eZ+/uY0ztK8pBQ1Rz6k6t2kz9kuUsvu6AQuNw04gs0vduBKE6MEu26qJXj/EIw
LtxZxvoUfUzbWx7MfFDfhnofkmKtcD/lJt3PabaClFait/0Dy/vCfaajBFahdSbD
sAisxELWrOdam6Eg1FxIC/QVnLM36KOFOsWq89PaSJgiHbrYakq4pZczFL/0qT9u
M7EoTB/Of4wMc4vNtiVDSXSjF9i4an8b6CIQ/VPHsBgeosmPabGt7yy+lXTkVt4p
BVM5DhnHGY2ItkrK5Kd1ZrYqnNMLvgRlPDY7+o3YWAPrwmQMZIL3RgpoM490ngzS
wA7/XyS2v14CYkNEOx4rwHeG/XLjD4IHD/n5jnjabcZxjaFpjTSIxA+UJN7VAxz3
tVovZnnTAF94HJyUKRIggnR/Y531BJsxLyAaEtMZrgokLT5HQxRz0+QllTt5mc8z
cle/n3X3+lSpNxlYJ7m3h90I/iHmTHXKGCQOs0CnOCg1UrCu8M+lb0z4NYXz9s2k
udLQlOw0GcbhbfDM6y1HfSA7YBy6WwGUwVJxzZ60hh6QAz0ardkzhUUV2WbZzjI2
YLEkkMEDyDujFDghOO3d6ttNITxzQqYOMKlSmBuRQrsaUFiHl6yaGs+/95G/Oiut
1XxWiF+nGwClJYYsxQf+mdzke8YEdJOtf/HSQ78Yn2nAwFpxuB1TAcFkcuPCnS6g
DT5/IFTfrMWdvk8fa+8ChHlApXoBy6cVxZsQpIcOYtf4hXMNcQwZ7VTpKg7ypUt8
oAyI4FQDAmuw1aR8NryCSDZRvj6ZPj7yIArgPsqkYYzz8J0r7loPPTLldAC7IR2t
sxrkRfmgC/XnC2c203YFTtPiD3+oTq9CHzCOxonn773RoB+dnsuW7D0SUecc8LL1
icFvkOVFYfLqd2lHtTlOPMWk41dvRc9+6SzU1V4//lymuQkR5k4/VMq6jmrHhrna
EX8AIkrEAJ66CoeJw1v7uIuSNpldbjEXgcGiWeWqPUu5MARyI2WWyV0Vx1+/QQe7
xtjZjubX5QBROOxMQQt7ZAKi3NQfGgaKPEtB7imskt4Fo3Zhyh1jB8Bi4GABEcpq
lya2brD9jIN1pGoKhgAQw+YAwrLhcFCNcGhikVKDCWZSzBQXeMi4RaD5ycAfV5Wz
YUMarnKjchtb4BFUS+B/wWBVVOeay7jjtEAqwB576zoc47cerV6m2L4xhgTjoO17
jVDu6f9snnTUSRPcyGLeGA==
//pragma protect end_data_block
//pragma protect digest_block
T94uxEPgdetU4m1+73LlTRusUCM=
//pragma protect end_digest_block
//pragma protect end_protected
