// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 01:23:51 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
trtQIwKS8ESKulbZE9WzDfZQcoyfEXSuakDcbr3zphz/s8R1BXboKUC5TB39ovwP
t4FPNmTEHADalof840Pw8A1tKDXzUsNf9QVQPtsCAgnfhsbYNfTF7IdDy14QXD1F
MvLRBTblf9hqvAjDUwioG9fBGaOc4bk7gmh+IYmVvso=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5184)
QKOrFU8gO77onbjpMTGZaFHUqIynlCNfyM/sihv9r1I+PK6OQOAnb0uUwpPpgnW+
zpijebKP2W6okZPa0vQBcUeZDcuUafzGP6yk8lQKf/eg3AMOzP3cktAsmdipJ7s0
+zjcOueDJ7CC+/sVq8/G2BpqLeB+78WOZm+Q0pvW1OqK+lCrJ4NSNcC0N0Y+XNXD
TJKbPnv4YfV/EZ+l0qOb441Gjw9c+l19GyfHQ8XqjIGnh7i5mm/RzIyPPPuuTFp7
x/8bRqAyG4hF/TSQRB53x5a5u8prFihLr9QVEgurChE3C9GBBczARiYMMUDIBtaZ
NfgrtvHDdnDGKrqrutu3cz4qFcyN0tXAXmG9Wys/v7ucw215MFlCkCQYeTIJmCfu
2OpqJPORBdxFuP/GUdFZPGvpdny1MxCa7npO++l0OuIVA+VCSelYapSQMfN2N4f3
9DzSGVv5wXzAlnDuSm/XwlB9x2JJMePWxs5DZZn8Eh5RxgOgZ/xqjL/J3now8QUF
/lZDX68Fk+QeQkRwNKLVszO6v2E7KFanzbR2Qnzg7tyVw/vX6qxcRuxSvPibaFUA
7pgBCc20prPY93Ds40/sxPLejr8pqTdqiQSCkVfLC69ChIOYO9FbupleSDz7kxk0
ITzmrDv28UguMryARvLFhU95qseop3l3uTjb5jarr3NTWkpjj0POsysse0zw2wOW
45g0o3Puhvbj6A8hlj0mat9pqR/BGWygodHNe2aTaFgTaznzMEVpn656AYB4fL0k
LhIpTgdL/7d4x4jOdHa0CFHPkQDN9fz8Lm1y4kIYunaT26VSHBYBse+nesRyC/HW
EfdQIBzgzJnhgLe9vpkARjgZPsxqK0nraARwySRpF1gCwUFqJ0JA7J7ok1xTL/hw
/4j9yZIYeSf3Up+aqclv2u/dp1P0yIJPUNTcqdNlOnqLGhjIng6QRRkhgH3sC6+P
qdMFYYBviOpc2l2cCOGtQ7SO3DaT2WRhY3cUcv8i81cytfemrkk0KEWdacYUf45t
U7EKgwfFRkv0CIvxWTJHGWQgkBWHqbD9RG7Ht+kh5ZMFaGiEm/4VGCJH0ieJ5rAv
LNMUYuplo5Wdic1j8g6oeLcmdrSTJilSdXzCw/SsOe4+R3dmmZohCEJSHHiRFMy+
abLz7S5KskDUORsZHHfMxel4Vnwitj1yfv/O0422o97wBpFd/1e6wQ+9SOkUqOyN
0ja68i3OcLPQLaPeT994RtI8SHCAxi2RK3ChE7RPwDfRXWaS+rHo1mwOErOl0JiQ
qywW41KMgHbtQM5cnFD5q8k0cYh8ynA8vc/Bbo0itrQohpuv0Le/UTpZdME8xatH
UgcSNMl/eZKdmxMuZRxk1YsTBHa8Zi0oQ5JZVCVGv7MaUs3dw2M+hy2yODik6Kqb
MstuNPwyqOUSlpsGQmYPw60QYva/pOQVomJa1AnIhpb94jaSIHy4+JNnpymjrFiR
4CttNODHnQZQFbvR9VHZTIA3XYV3KzbgwXNMMVpbnWsoNTOy8T8PwwVINvwFKwS1
815wMyRCQhTlPBgkjL4ZLFsw86u6feO4E8fZY5xmOKZps/mAtPo8O4KFIMurdsgT
1cE7QYeMOgT7ZqTCVLer+KH876D+asL6B1xNeY1aoFIf6Zz4+cbNUPB72/AGAKWf
ArHhyb8+nMQ6j0ZHptz/W0H95eB5aZtehRUtMo1eMpdpYgg8LG289yB1oO/r5YC5
CrsDruCKvOQ+U82ICG1E6uM+ofWlauGqAu135o3TQ7rdhFMM6Xs4QfQx+fXFFRJC
rxw/4LTOciWWpVeJTUjANRCzMje9uri7i+JGvkjnvjIMUpf/0Fgl9M2lSzluD1HH
LWwkuDvzuQUyIprz8nl8K7XsLnqeX8bxLIcjhf/nOoZRnBTPTH8jBAcduqECLFXE
oA8CvKn0kAHHGxnFV3Z3glaS+nZxVTZaO1wM2Pho3I/57OcwhhiAQCJcR0saoaAX
gJmEnhc+lIeTNPEU6xz77ZsogvvOkGyT2hzqREEmHM+rt0AADX8SURf5JS4rLAcS
6rLek+k0RCIzCySSfMlIfe6BVclOw4bMplCltTz9O2gS/HNRQ8NHHGwFMUovJvMq
dCH/ZW+YEvPk9B8u0xC6C70oSl2hrQnXjdLfXxKfY83sOB3WP2uspU94brQZP/zT
ZA0up5rU6J1januuwTz2lqc+2jrDpGyGQqU80Mmw5kmTDnGXjg8AG73ZH4KTsvb0
Fq0T89ELzFw5rY7VfmPJBh9mNujcVZ2v6L32AQ8DdzWkueCtjnvgFdRKUjruLckO
AySSvISEsnkqi3WrhsAT1Ghqi8YxbBWs4qJgXm/hTrmHVPHGsySim+Kr71kUGrP1
YyWyikmpn2ImqPnt+NxfoiMjmd+cqZ+IrYiW1IGZPUHlGUPXH2dk3OHRyu1qzm63
d0Ufzs0c2m4awRSrirT2mZqjgCoLS4iTf5SS8MjTxqZxnmjXAjPvEKZH4+oVyQc+
BjgPDSG3Vdb+fEb7cG3E1+CVmm+gPEoak4D5KcqW2u8OKcGpsdZqu3/AUYXjH7BX
ag3S9MItgteIiL/TKQIKybLQPpH9TU3cvIp4IzMlVIl7pEjq4gQI/YOiGkal9rIv
mCo6va8AMdfaf7ctiuJBw1aBuYJeaBuQpXbH+JfQ1ONAlfuE22x9fVu5cfPyefqM
fSv09FvDDsgSI0SAHBiM+gODZuR4tBeP8oxD1vqSTt60n6z+U2LesudU28vZOKv7
1j97eZLQhadbcvFqiNdQM+IWkJ//cQTFWd4Cc5S1moCa+LjU2+tqSjl1UKG5BDhk
crxEIGrcUE8oMSTOr1filmwnF66vqwKgNur+Shld/ZRBybdG8MBfACPbJUXOqund
NYxZqp3CNgh1Ml6k7sey3ULOEFMcRBkIyCX0l4sWIOnXDs2l1lOlNql4f4vdfzjh
WmTIWO6hBkxgMsgDoGfFSsd1YNQ8WwwDyIe+rtQID9e+VznaXlRqDMN19R7qpV3H
uk7iCQM3VzQAk0weEgvE9yyEMJFTWFfGkzoqkNo/Pss/BLlLSo87xBzuu5oLRBj9
z0s2kDUyRK5ogNLkDzbM3+1hMKCDNX0JHOnCFR3UkHHbdY5cpz5MzoQnfRIOHpDW
a8fEYftUfJCqsASX/ibIitGCLz/uRxOnpbq0OxZWo/1O2ptLRTMfKTFtvaYypBOv
j6UIkhowXCNLZtkCV87lNg+0ZTswGw3Vdx8g3ilaAFwaN0eVhJ6voLz3pQHNyAKe
N460LLf2ShHYSXQcKwyUxpta8hBqsHU818kZoKfi8LTVjHVlhf4kMI/C/A9tae/S
SvYJk4ou33I3uDN1QIQX/ZlzmMgsSyHDDfMkeFpN1aqr/g2T4wrIQblZassU0Sxu
phPUfCtdCGe7VfTWgJLiFfrAqeocP58t80ENybGnHnZ+doacVyW47PP+Oi/UUTtv
UQKec22dUTlLEZhEO+DVW/Czaxshb5kPDYmivMhIVJFjoxt/I4R0mDhEfCbUxXmX
JX0yol+bu11z6UtNZPg7JRjPxT2HoJGe7m2CHyPWVPdIJD+YZubpV7fN/LLt8RWh
ruSQjJxhkXEWuOXZy6h0M/qgZK8RRsemrgJsRPsHJoO5B8YYjqcJmc76m/HPBcbN
HgwufkWatuGKskat5boi3WbQJKY/jHqtFDC9P7jiklYaYr87c3SZP7Zv8qXLAVC2
6oC8ExTsc2gyb1tODccWH3T0i2tvKu3yOJWTvorDsUQrhFvh9L5je6hEIPwrEoKe
t/YBs4gHLHN3ODraVmBuPuOvu9Ayuv8ZDXl6yqIASd//8/trc5M8P2U2OmU4LWzX
LUKVrxW7NaXUtw63zEqsoQxxCQ9mkFsaanm+Rf9TnAUaLEznKgDQIbLMqQapzZ/J
f4h3sFL3vUi28849HVJBjHxw3FzgYoXhmUjtWZuFS9/fvpblKby3AAg/tiVxo4ox
WR528jWnWZw5A7fn81sj3sbENS3W7TtLjwLf+gRq8gYYxWQmoxKlJa/QPD2zuYGC
HPSDMzdQXGNsZesJ/Uy9hkWXUZ+D66AAYlHXw/Vq3zgLrpBGnIQh1Hqmexl27ikE
0KhwYG3YHcyZYYV+WW9mM/ycGGKa+NJovrOLASMX/Xk4SMAQYQCKj4kcoMQAK9u7
OI9Xtt/NdM82OG7ZP0PDxcPs9bPrKS+nyzKmCtAiy4e+jtpT8dWGzQdTHW0GYy7Y
t71VHBnDizXNViauo/J6utmUVYMm8oI+aalSNrTxIrcM1I8nvZxKFd3DDVAe4qG/
onvm5POfFdB9BQ5WTeVthbXvPD/V/hEZaB4dJsHtkhKoGwxFSRhFMc98xd9EWupk
ZrIqT9Ln1bHNEaVU3aGl4tqoqNRmH03dqQYk9MkHDM5Ywnlwr7MaIgwd/AdXt8Wu
V3fMLkXx2BSeO1pZEN+NBc94HIjlt0+TpvzeWqXIDZTiU5Md/ZVXGcMViSiQwZXs
EUby/N7/eAxPdqotTSl8nS3w6zB8JyRT1w4Rk13QJ+iYDHtcvwViP9VTiA4XUqYu
4IJdA/SCArrdvMqd5tvawl246zWOTDRTcFzWk/B+ddSLbXC2I72Vl46cz6mcupKj
1DYCgQhOckpZhNYwYW+Mm7y6N6n7RkB1EM/1d+sltKePztan+QFTb3ixptt5hTDu
rDCQlckQUG8kF0tPocQQsTqbcoV6EmmJPRUNZIsTeZX5c/2mKbSTV4ph+o/vQTkQ
GYukx87HdUPDxNL4w7beKdhQMVoxg//Un6Ki/xwNHzteE+shlkZQgMbLTuNji2aT
veKwwnRLRdv1yJttjGn7akZKgIttT3QWxd0KmFi7ZpF/GsZyqOByS4UNcn5MjKsl
dAdJVpASV3XiY7wb4bpq0+86159/c0MsvNtXzokZh79qPrbkNmmftOGCnmp5yfQx
NoLdOWeGzscYicnr9X5qAk5v970N++zeqYbmhrqWGM1Uis9KW76R1s2uC1sVRm/L
9WtUaqz7HlxYkO9gsS5V0kvlQRsbZQDZoWI4K7cSaXmJn7gOu5ZT9KAg7VqnHXWt
XvlZ56U9q/iywz54VSKG/m1tLu08INbK1SaGq5DJLPSN8roToRj91Bs1L/j49Nln
bNdLviaeq2ZwjJJ/JUhmnzC+BAmlGPkrQR6OlP+P/d2cbYtrQZB+VNgg1smdWnwS
xXb6Q+TM2M7mtBEHYpLMrAKdl/NnuK+7bS50XkbPZdCvpJa1GxzTfgGFdIORNlE+
gtWMc2SLgKK0toqlMLo4Wo+sHsrHpGaVFkpqFMZcNdhsWz2ALi4M2MoRcUdFHoqE
0jGXHd/baGsOAZ/y5S6oLYkdxnSAiBykK/1vGPETyllkEgGjq35JNVXL6sWGrdMn
+xAAsjWCrnVIRTjAfSXLr3QCTMqLY5bq15qtrzsANObO0ZYVhVFATd5RDQzkFv6y
7NKofoC2uj7ADuPvpwVOaHvKylm1tdz/FxRuJpo0zNnLUUjGVKLv0RlVi3pg7uhB
vE36pBtyGRK1f0O7y2ahD94D/BBAEH33hkkvKWqETDZIBQ7eCQ+D5Dh5MKLASmWr
dlEYO1xhUmoEpP1CYM1oyehMxhbCflx0EceOY2Q3F6FWppoQhF968Zrltx4LLL+M
6GOiqQZwhAmlSHOvEA7b7CUanUFRxytcXM+UNbIRypi6oSVMIztf1gN/Yyo5g6V3
MGMBEJwx3Uo5lspagtmvG2Ukg6FskR03KhkY/8LE1W3KGC0oy7rXD4qtIytfRK5e
681UMiR17IMmganJL7XJaKSSGzw/UAZUZzZCW4CmKVdgVMsUPEuXE/6B5D8D1hYl
xOxXi4B9ycoIKrWAPUnPmjj6daESoEQln7C4zbonDG9CKXLtJUF6+hb+cFgsP9EA
HK8AoWXgHP2KnSc7FFD9cNYU3VVGQkm03t5IBsGNclwoawN1sXYF6NjeDNjZPIKm
H7pzP5c7A1LIqN2lbYFYFe4j7Jdr/x49yDFGWA5H4TW4jalbpF1wGoFPmNPKX+b5
7OltXyQOzJ0PeAonCI6nooGf8czVLHVWrFoJZFVehznrwYh0tRJCi15VOkuVeC4/
ED9NYjfxn5NDoHLl60gRgFlrqHhhUKuW+3aEukepJZOrjsVIJP+VF4UOSes3nPo3
5rcQqZQhpX5Xiqhu1fdrLDaP0QBj12rt4EL+gBcvzYnxG2uhlH5s7wu8CMbnrCxE
PgrewuHT7dybkcNxbf1xD1jFkyYtl8P11jVE1+rIu0+yTFRirNSuZqqyF1YXCZD6
4/dc5Aw/P9QvHwz+LTH51+xnpu1fTlHEkZiCrzMEwuSCPDgZHMgV7BoBevml2z5W
wXo7T/9FTnylV1QK4xGSR6JckZClrLR0wlkzpyXsJ5IjnEl4WJaWI4NoAqEzixCz
q9Tx+0+k50x1IKEGO1WO+pHyCaUhf98slvFxGDbA4NicdVCvKchtS4942Jp7qdXl
j8peAP7S5qo5jOccHVo0HP551QWfPR2EZ4Wp/SP932KGKCaDEx6F5DbTRZw9rS+P
eXcf/gqGgjIsotOa5S4h6uloL9QHb5bJJEGTK0yqjJqiIpPf6DWw1NBaDzxR3K77
YxnpU9i3XuzzCLou4fyCx6M7X02xnj9sEoJ882Tlne9q4FelCYu0aQhhFJ3Er5dK
8z2eJeKrkNzVhC6u4/pXUlwomCQyb3sOgBKY3M1DxV4w86GyjEtlKV6IVesYggQ0
H70UoyUAN9/XVGK/vuytyUKI8Fp89Idew9nlfVMvK/UVh86GM37vFmfb0Iv0Oy8K
MWLqJww4nJc0yYMABbYX9pjJlbh9crrQpxKeMQrqmA8tBAsd33UDeslpuTi69t2m
DoZ6304MQk/uq4ckjadDtwwAVSoznF2Yd1Ao7FcdzHqR3kk+Ikm63vHM92NpsDkq
`pragma protect end_protected
