// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OVvvYbKsbXbtxZGXrDvdAu60H5H4dx6EJkw4ygP6/seMf70txxuw35AlfT15Zba6
GYtTcmZOTujEkV8nADO4NdOHT9Utip9ZbqNhWotK9G9uFU358melknom4Pz4nAe7
bM5UPTPm/EkxnEfNzzFDBEpQv6+uuaBwguC9t6oSf+c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5184)
E3VuGQcS0qGpB2j4mIbBKx7ZNCIlHO/iHCZFDswAxQN/5jml8Go11YihTkwtNZB7
yQ5cuXTReCxykjV8ttUABRgG07cgxOR43yEOe9iNCOsQx79HqLr9xtn4ETlvnmQN
hZRTauPUcHxTWc+KsO5fuF6QKJaxjIGBEIMN4PRqEbQU/3CwQ8Og63ppGvaVpK1i
iBRhLsyDWa+H0D5ZxzAvrynIdyhA03Ws+ezEmOPY++s/HBMWSwkAJAefPBufHC4n
80pL0tygf0Me/EIYPOxdmvPa30GifWxItv5MS4hf7NT6iZe/tORSgmz+Lpl5TLVb
BkC5ZuhCZuEKNgnmO0kC+A7eTviTS7LH7M6bTkDK8dLSqy6TP3wExj2QcJd9sXfg
Bej/ROH4dsA/aYPVUG3YmHkWQOzczalPRm/u/zNwATJ/jmw7EB9SmuflvdDPuLTN
d1r+BwfvdxLHyAjHVL4T2fAFRjCpC56eAX4QlozzxYMTSNn4xKPs/UCM5x4snkbO
NBj1cXEPnIHNbmbKD9EYXZBOsp2jmgMfsK5V98PL9efT5A8Dycg+evxUZjJihIpt
QGky99FT+apCe+5zysb0VHglyeYfR0iJLsRVW2abUfUqWOst2OQAEibuyZP3W+4a
E/xOtI6zvMGsYJTbnQAxS+JYDotMU7lLxTHC69wZYc6uZFjofTGq4vzqUAC2dWg2
iElaSE77g23f08PVcRPFickz8n0ij4kJgKasP7q8B4ApXTeBndUUXsP+71EF53IK
dYoEmrIDIfthEbmVNpF1SnOKxa+h3RREgojz6sCPGju9cVmuDuPYvqoxFm2Hd3EK
gFDeWUkcfGUyDw+TUauZlsKbRJunXRusczcXvfZ78XqR4Rx1ibZZpzv/8aUQ6CnX
THHJ9ZahkMvAJ+Jp4UwD7kRcOf4IHk3OxeUbIriXIgVirmRxW88PmkVSRbEfkqwk
jTvLNrqZg//X16kOZxX1GLA5am2aEAgWyN67pN3l9E8kT62JnzjJ66Slm9+iYTcF
dUdyoeQ6jV3Zn+lCQ4p0g/e+xyAERyVDeSkzeWy+J+TkZMESdJW63P3AeoNtXc7/
SNt8ld5UknBatyQHsHclrTc0l6KBkm6zd6lC32bcY5q+U8JkZ0x98MBJiDu8pNDo
CbPTW2X+0beaoQ42LeQ1vMYmrdJNuD/1akrrYAsSXAyKl/8iRa68kIWOBJhApVLh
GDtBexNDWWbVhv2TdhHKJstrbpPjXAHCp+4er1OH+/zN3aBg23bLC2sqW+c4MN5l
JMRWpbxOO8Uixy9fEBmeggu5KuHq5kitwDiHmNK06Xq+PDOWhubJeSAJa6BQYk0/
XT5X0EfyH4E8MXoHtFEHfKgXChvYmTJbED5zlYA4F28r2sk+KLIwFqP4lYu5w2nH
GevOsApk5HkYWVVCFKFTXybbVQGZmyoZRwBceQeZ5FGLMmrA+it38sLCn4Rln5vS
22XMTVuEDZlVL/KDHFR7eTOyOXcCx+ItOyTaPQD9G10QPpxcprdWCCIEjvHx2MFQ
Qhsdg6CxuRohW3ELM3Sru83u70rT2bS3fsZuUdIp7CpDq/YufH/Urb1DyPY1w1H+
fCc6QbxXEv2duYS+rRSPRr+j0gYj4/yYSNQzuRuAYXU8QUx1bHaAU5vEdGk61Cti
10ZGLiBP7pT8W9VSSfDLxPt1FTYuXhZ1xxSwm3aCt6ZHWrEcJC/fvWWxjEQG9Iaz
OiClmfFPmZWTSQzCJSuLXhq98cVcn3L5EyBd427KE42u0VxyxE1fi9zolME84j/A
quIJGQILMICcoVtsExQy1fICGhANdJYXmCHZKvYuIlkyM1Pzw1roXO7ZgQSiGDur
mkps6zjQES/asC5eWi7xaqzdsUCvvBEvkkDvJMwkBeVRIwJ4+gENqoyYrUykDrMn
Gv/iXXRZenfohA+W01qZ2EYp4gOtjz04OewPTjvWKFhdqgygxxXraB5puMzbvZVE
SEqCBSdvYl7sAAxppz22/I2MV24M+ok16iNrdTqWKidu30wWLLRV1ybZhV64epU2
GDXAlsBX+AN9Ifu4fHFRRJbUY94fEYUPPGIvtbpYqGVQKtls/vTL8XSRdaXpv/Xv
4h26E8WnoTcIC+i75oYuKR4azUAwT7m8la+oh9SXDDzxi7EHd83Za4hPL3+jN0vX
S3pm8Wkp5V0yypUzGZEK9+ZDqmOI01LwBqIdxy5Yxe/zbvoZGrTdHiYAjE3CXfZb
XYFoE5FGe8bKtzHhwDbPbLkOSlDtmAGk6/nXSWT/4uyJKUZlVHK1u+Oaiaxh76VC
hpp86xjQrUdNTzPA4YCBPt8VqwsJQqRJ9OPnr7iSPFCQqj0bdpG3PlJmFCwa2pPH
e+RipxxdxNwd2INoATRo9VHEkAulP/XMVAcUTuhUJs8Jf9/onpqDo7oXSH2wprfK
RbzvesfWPPVt5sVWsHsG2fce1vPJmScMr80oOmYAUw6dxlViqZJehvmPkDaNE9GC
yRqcJgn49YkpNdBXtFQlW3JENKtWT6Sd79YXRKYm4hsPGEQCq9XodmML4pRCmJv+
iggdDQ5zLVAxrU1Czxq/qWyodD9Oz7Vp9k6ypN1RSYjx7ZpKD4dE7uTtlOFCt7Zn
wAg6hwJvg8fILw+dw4G0eCBhXMmq/1SmiT/5RYbaDbcOwsBbn3bTXb4v0yCPtFU7
YlRSI6PV+Cd1HMQx2OUitqVGqaksbqrJ5+mHllUlefPPmVUYnke+Ua7PvdpvUPPL
mE6j620K2W1UXZ27jmjMkWivW0adma3BE+0fZBgxiGqy6hWKPaJBaBBXk/W2nTF2
j/UcO1euBafz3LUZyD7Upz2jUe9Waqra5HKx0sKDkSNrM8G1caa+kBc7FEIwbaSC
wEezMPWbhuikCiiwnGcU3Wre4vDDU9VUYe/lraMfrVyFJB2NJugG0mxogERotHuG
s/pJ6d0pXHNXuUSmf40gc5IV/7iBye6eVI5k4hHSqMXHx2bMWfTXq9Nxue9ILvlo
AT65o3n9aKSa5VD3Z9eZ8er6G08SJ26CZ73Zz9gJA4PZU8MuV0vpTft5uPhR40jH
kUi1T/0lw20o2ZT0F64WSzNh/pAypzuxI0SeY2nuFzwtjGS5SZWZjIeZox6cQLbV
3nVYe+BEY9QumMLBcyxnTQjdFW9ODIqGDFy+DmiIJ/DldzAxUhqHpZQdaV45WWlm
7E9R+djLw7b8HCza62FDJ+Yx8M0+4Tu5N3de1Y57otH2LW70ZkgV6psHMR9l8tyW
/8qpVehIwSUHRCRx+3fFTyiJ7S02PIUql0fsIi5s8PjMhZNlwtOEuMfzsEyjEfN3
bta4/XXDQbRpWpLp3Z82MTaG+QGzjy6q8l7szvz07Drz4SddheUbc/vMX8x6+yyR
oE9tnm+9gA0PfGiybB0SUjW4EfECjw7gsyHMs3L9mf6PL0AQn1HGdxHZJ1XGqhlv
HiVPxPQlwPRXasKtxJZ+v7zNjkmKzRZrb1CJnfl4iVaDdXBSIZ2J0kw879B71Bqq
RWHkQgAOo8cjxJ1roHHyObAr4HJCFRipWujZ3HaixHzwBaeJEc4uu90U4nNXsFFq
M5k8iB3bnOiWQXjXTf3FJHBsacsoa+tzdnLa0s6ed1xRVJHhtMcEgDNHW4FzVnD2
WYfwlaZC4qOEjiOFFKXIP+op0FaJkOjniL0af9WSVNPMWAy3tTFpDQoS8txIOTh9
Gs6pfPR7C0I6gSCHnEqYQkmyiMQZWvs3ps35smBBVBPQHVs20YbaQr9SnjNcfXDW
E402jEGTc2TZOgaF3wd1Vkeq9HogL0q6gABPnzcz2IZY6xm1NirEFoyPlXhjGvgJ
rYj7QwkqHNHZhAcp6SdDjFYYk4mu0O0Ff5DfJcObB4jcY67ciI7CvJNem4fG2gB4
iT6ixgu5NcMF5j6uwrvplKGc9JemGQ//VTVJKbJfoYxIHXKfjzdW/Y8HqeUv7hRu
nh4Lbd0a2+VRDUvGCjUmLoHUgd2ffq+uy5cXrMtTXw5grZrZgarYXExCPokkSDGP
RbPperQaOIDfQ2nQc9lpg8FOQ9Z5Ttcwrr3MIGV9CUaQfzRlpZBQkX/WOZjhmzuS
6+9nP9Dwczm68KlO1bzVTNBpERPuHBzlf/oxgVIlnvh6Cr57zrlHpzkOaUhmWM+4
gNq+ewZUeQHWoS/cVEiHd3koSOsHkETlxvk52cO2cnIvduTlJwIt9iER8VHk78bg
2ooVl++Kpq2TCKVnWrJBgiST3MztN6QkwC8vTPWpgnSD2Ti2uwbZrtXfd9jgrxl8
gsE3HaRmWoZMeG2tnn7h80DGh+07wDWtdBc/ozFeDf5IPWmJqn++MJtZpi52Og5M
o8CPNV32Ww7qv/MGLoK76jxwPfu4gWFKU7rweuk0SgPzK31j8U2jwD73ptCs4Fz2
/JVbpA7TSALrBG14CHkFFq2UTD2UHZ5M0PnD5Efj5zgMozsjEb0m8hC86qIzY3OJ
pxXl5Kjc/XWb16qRFT0FWCCzjg/d8r+0+fCbpSS5CedVRmB/NbU1R9TL5mtDwQww
iO9R9sbJYMadaHHEvUW+1F31AocRuj8mZBwWhJDthQY8XpKPa/xoVP41NYtAN/Z+
/Yj1Wj975hLktzHBGcUNIiSTV9bhKJhtJG+ZROKBjYpasJjEuxev9Y1mSsHP7eRk
cABoWHKhuU7KWT+VYA3JbaGckP3hNk0bT0oupbdEHdkmdBGiKVCUYobZVUtqOi/q
A3725uo19Kry94nyolWjFtlO0rsujjdWzjFx6j8VGZ3FfUEgxUKD6gx9BsbhlzMp
RjtOTuN/SapsbSPvMp9jBx7nj1CRxAVwm7xgae2IQqPZ8TGpD4bJfh6tKHi6W2Fj
/Uuj0r2v1RjqAra4T6Go52fdxr+NdkdxPHfEhpGxX76jGZFhgdF1UhHmADLoxXZm
6JAmMyu3gmN3qCe+Gj70aTsJ/1pgA0Mx7A017xCyjCVQFWM3X2US0W3ikcKajfpF
GLLOt9jbP3ndiUdPhmZjdPoQBJ78GJ0QNab6qYgNTwhuozUp2jJVkI6RFX2/Phhs
Dh7lBnlPZXqmDoSpxCS7o1LnZcaWkLjJfLgRNqqil9IqU1qHjACbzrmkjs0GwkNy
fHyBO9HGxAuROY1yes37L2uZmFd9Dynl0rmoBrbFcYGdw52PULea+g+tsO4FyyxA
+QatQO7Tryhgxg8PFoqGMmS/jB7gLqUhUxAjpHBhPEAzhpQ5smMU0AdbXg0RoDZL
IaYAvhwYF4M+HQY7csvpZelDC7si/5ftTzxQbiO+3O+2I37o1IsnjScL4Gveh6dH
u8yRJ74tSke6cnNBVLf5qrj71fGekxxLSe/3kLs95ZG1gjrryPg7ENjVCOAXjV9o
KOJz5pAt4zZW6tnjapM0cgikIRYJ2/1EtibJA3D8/Cj0EdrcGRNIDF1PBhj32xmV
+/4Fl8wfeBTxzIy/h/RF5v5VmvsOY/X1u94NeNEm0nYQmIJhE5fjeUdtmgMgdG7u
O+3d7gOVv5bm1YaXDEku602OgEonrzyjvwHsRl6WUzxRYZsFP/B5FXhIHx4BB5GG
iYHUkys3FGT6czvHcoQMZ7elEYMPna+NxOnvRPmmRHrNbHBjfwR9X8v2xMw5FNPx
MEDqffYFW4fn+0Swxm0kop2saMuXPG6rQEHkxk5fD4FMi8hcq9LwldFLvMHP4wcc
5KXvxPcn/dH0FIhpvrsge0FRG9dKFWgvR48R5BeByzbW9f9389dV9qtqb5oHQzd7
ZsB459brwMZYR+L+JQDwghGm9HZepKV/eGLo93sEEVaEshtZ7fBHnAXWjzMgWKTK
I3dIk68U6WmaU9a20DzKPFko3IseFpAKcMXlvq810UKFNuQ/3XjCQGKlZb3kjhgs
WiWTzy/0Pgk3HsW8OTOdc6m4YzVW5ckEUpivwex767ZAOp674qB4huUktoI0g71O
6AhZ1hFdUAi1yjidJpDiP+nBa3NCDVqMHf0net+DgYD9hrWStniDPNkC9/tcClDu
dx8rTteictxnFysFABB4+1r/bHRfTZU43Yp1PpH2t08larTMbF49pC5y15gmvYmw
otx3boPjHQ+zi/S2TS26cADP50NP3ZiM47C2dLLQT6gVq+Vpf6S0OQN6huacjhsB
SEodeXh8RaeM/nU6UbfTlJKJv9AJvKSIJpdcDe0Ca/wtZUL24Cdn8AQo+BDI/v5V
TCxDDF53hMLqvlyVA2NP36jVqsnMjdZc25Jd6abmtxMIxvzR8FsV9P7r0I+0VUf0
3IY7T/8QV5NKUeaIEFGYBRj9LS9ldQvudIEl8GIv4hGHwDttgTVXZm6R92aLLNA3
Ekrd7qrOim+zBoBPyUse2m61X1O4EhVyiEmfiNwKvsdJo0hlrDqB2pqAvKmT5YkN
4FPp+C3p1GgB1RiNeSCT5MJrtsMMw6kW9iMEYsvlUH2CqFOG0wP8U1O8tBMe6cJN
bUFgCa1yXhSq/5etktUWJ507beVZKw+kwzCYdrEJRZMFfjkY5lXBZqqJUkjX4hnr
92UvE1i5YA1MlPOdtlAheeHs9AsiqG5oJ30C1aY3mQpJ+tef0oiKFBl0lCjXFhFA
66K8Oso25A1gGfcGS/jhYcl7B5g+vaVLx0c+j8TleLOfjiE2cS9DcCOFDuM5mzVm
nAC8ke2p53eyWp/zf+1N7NtvPMpRNxq0FfeQtFoc3ULL8xFWqEMrMPN6gce/emt6
lBTRJDAfnif1MPUBBSV+S7ROqtO+ozKRAND4HNbKk13hFmv62wEbQI3G9OT7bFIn
Y90yYZIISq1mPJ5gs2VYSEcGPT3zxGAdjLbhJ88bjYBKqinpnZXhtWfqNy4JyPeo
IlICAKxfd6kHUC0VHC9rm6uBlLbZTORl8D37wFcX2RpoFgJ34Itl28rNpk2/8Vl/
`pragma protect end_protected
