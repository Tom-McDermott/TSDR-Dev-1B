// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U2SJUjnPUznV+SdF+CCSKH32kUyfYaE9+MCQfAIPL3KrTQW5S9ZtZtzKSI3R4pee
FZog1MEszB0eP7hkkJyV24yAa1fiJkppkEjDP2Wty7FeBhL1NCCuGhOhq4WJrlNp
vmb2rXgKyPaTNsB5g/dTtP1FBzaHOmEsc1nEbkmaHh8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6464)
dKiLmkcmDMK2KWedzhShcgap4nHI1BM8AYbEskmyCt7laJ/8efyeBEY3OamTsP2w
UB2NKIhexL3Fiqa2ETYai5+TnGgrJKJjA//AT3/loD1OBRxgL1JjxqrDahd+O9TV
Zhd8WchNyF23vvcBpox2ZBuHo8hJIibrPiY34XMXS3GpkmnZtnbeh0qg0SHZlfIK
rEqOgwUwiUl6bdDMt5xs/KcPdizDW6bP6gbESmJBZqkPwf3XZDIstWs1ot1VMGqt
vVBoIax4kgW17m0BxAgb8RBEaU5V/8IHrXL4JujZrySLqN6we0FrJKlP1EsPH2zu
Pb5H0AYXbGMA0S4ZWRzgge9lB6VUInvkTG39MuEKGme72FFaZHcaP1+MYaAvkmnl
63YPPDixFITvCs73bWK6xe9fHa7e0lWySLP6L8dmmHWR/fHGeDX1vvN5I1GrRQSY
0lJwyr7N6BIT6W9h1YMFKlD8ip52rIvPZGoHdjng8GmB9+9aFAa9Mg9oWAsguSq8
CHr955I8HnR1gKOLqvD2FZmyox6X0bABIfob/ptTPEbZpBe51D7SgSK6rKVarorm
n0eHfh2hurXmFXBsy1Uwf+4zcGgKhtKgj6InO/goY3tMGeioYbCBisVDLlOCk0IC
qK3rqzhBGzGt+OETpNk2I4CXKUF0+ajvhrSfez9Ww6BknDTLiwwgqxJiPktU+xo+
s5LuJpz+bM46gPV3bZYOybIBox7E0o9Lp4XfrW6MP0RadNEy1ieMuowIMedXgRVS
pB2qOmpzZ2LeZ3lBkdpt9JX3lXNlVWKutDa7BYK+wjTLo8NB30KrqcPd9vWdFHw/
A2GFST6TCon88z0v3wMws799L0WR02C3MQSIPczQlvvvo83dcpPBWsvjAsicSwwU
7dWXYCGt2GfNK6GppdPUr6m76gRNTxcDDV0oBdvVeHTLmhA0sg8HL885PYIBMvUu
yuEjd58DOJfyVSMMRkbC2nwiczi62WoqlLzThF48D0NrrK5yHEGONVV/YMDiaXef
1eOriy9ufWWXdts1BgvS83R2/arDMwJWfmcwbN7EYGHL+GGd/CwMNz2rt1LMcTm6
6jlH66smg6bN1C9C8DLGbxr+IuzCJpAX+vsnSPA8KyaaQWsJGPtCU5ti1HFsNzeA
cHOevSxyRnNNgflp3HYlqBVj1rVCmFbfBBwr3g+GDr5JVyY7hu+b1XjSEAV7LPL2
aSzdClWEfvGTXyO8IAhqFoYLDP2FTBvnQUf0cZHv5MDDoBPMfYNOu2CLOaucqcls
4PKR8HG4pYygtr6txeNJOWv/3zx1uWuMbutqQ+eYLgJ3VSPVk02QsE71zn8hJ47m
negxi3ZozTt/xRQ+HNzxQt1iuBME3Q9wpmG2OCgjTtnTrHzjFKz4ef1j6ZqZrM83
aUqXsehrHrwWpIA5twCL5zkaDQtXlOFD4C0BriKIHDMil8zFimzdFxocTyN8yj35
w1+UQF3XAl/lJIcdEgdt+iCX0JYivGVRjpIZJcdawtVfkY1nBidSwG6ZZx1HU3CO
tWB2m39DW/gfTaKmXqiGmeXjr1DpMg2vJi5Dj5pWgTAmbeD69ypnZIIWHpUgvuPJ
M3niHG3czGcxelMtKfQGmn+3NMl6dw0/XSumjbZkBRL/664U3FnBi8FDJkgxfK8S
Bi8TFJlufGCS9GGaUEqR2kIET+cR7yvbCAz46/4n2JW6S3HK3gzWUckeohiremPv
x27QmbmLNDebYX5Un7ETCNXad3J/5kTc6nkJI/+4Pw89+bUWx6p7vBzkK8RzKjDB
84X/FPQOBGSsXdvmxWXBwFuAVvxm5PVVqb5ucV1ZTt6KRcsF76AXMp6B4gtOpfd7
yyiWMVoS5+XaPLhlhZKN4J4huJBKZ4hnklXoe6cI0ZKNQM8r2NKDdmuInvE6gTfR
0uxjJkmjwR2g8EhQGZzHTbPJzimAB8F+yJmKqNNSujz8tsgc5TZRqb437YHbhlK0
/UAvIDiEmaOzGhVhlFhGVeOeLfHv2EVr5pj9D9YJ+dkeaKy/l69hFsAHWXYdULWT
vlyD4PYDvZJjWZIqIbty/OcndHC+k1aU9uhTUrmOP8W9wYKBZ0JlE6eze3l87qbQ
HDRifChz9ewr5HWfV88WfRDS0P/vE/hR0ifsRVcKHVtbdw8oQRrzf2a06g0gTfAC
EtydsIXHj4QcTzz/++3bcxEGccLYJPBHQ24PcidstiRJIh00yQZS7ytBCWkKy7qb
omSbRdMtdarS6sI9e5bN/3k+n5ZOFOZe5nNPdXz5X81wzm56QdoOVJ3aFpcL1vER
nFMZikfasXsGp63+/7ogDIU4BlMEl2X8cEDtzkieGqa51KPqhIksB+JD3Xhn/TCl
vahNN/J18o7c/sLfd8Pop6Vxuoy1HkvJiRSgzex310vsyIerRNKrJz0DPCGMhjl0
f7RI9okXZicIHif0je3Ht0m+xV778piFeZEXtjm9FjSxXj4f7G11dmVw1E1WZMeF
s21lj4R5e5dBlrL6fmp3oxSCQfNB92ZsxvnVH/I3pMuMH2NJcBBRS85IFXAqlJkF
tNpC2Ueboo0f6P07rDF/MvkhVqogYFNY2btMzg95AACT434hSwoONfvl5Qa0REbw
RExTlfrDyLSX53iaRCMAaCs0nkXUpWSGFRlppcml4dYicv5w1qkAvrlNyHh4LLLh
qqupQqCfTbMkd3O56gI8AwM8Ljy3fKL8jspZ0tGarFdEUrGehRrmmvtuOiSyD9Kd
b4prWaLcxR2aAGATgWYiUwK+vG0ZGWOa4uhzte2CBLiWwIzUKXRJWVOYijDwIUjj
b8+gSNGxNm7OD/FYAx23FsAd15HFgvqK6KsevGnOB4kddHHV0nW3MgVCuUMDkZeI
gFSkBP1sBk4eZ+/+Wijux41sabwtHLFEB/wNLms9wntS6mL/TIaQtZxxCERIb7o+
eCqpCJSLmuZPpEkGvRWGeWEn0ZK6lhlAl1XAucaypcZedAj4ZhW3ypx8Mel4KP0e
9CeROry5D+lanmA1T+E4pefuLLvIwGzWzTFwvikoQB79rjuYMh1QeZ8Q2VdX6T9B
3J1dAlIlO9Fu52PqMxuNCpFnikDjSFOCCt8tw7Uy5UyE55v7l3kOjzAuJNJO91Y+
xzPDw1jdBQHTqhGNa+d9i/CSZOVZNGYzBTrG8Q14X6POilpgC1hioly/D8qqAk5L
1HSSWr1RAxt7DRHk+IfFPg4RmX+FSZK/liAeG1omwDTm/P4kMiLnGXcF53AWFJqT
lDjb4xgFuc7zkRH3mtsMfr8cHoPkUTg2hH42YmVj3/RW19GMTDETG2wdAf2rM0WW
+zYT0ws04O38s68HReRKVJaiyLGl6G3uiYiL2Aj05LBYNKnjetHKAxKsW4IOMJs8
Rt1GH+VvyjZMyHxVcGRtbxtTgYGg7fDotwa5u2yJBaISkoq74B+D3idxwVEAsRnI
bfrVgsXxcJuzSlRLy0wbbJHgpxkKxd+Tu/coHxymnpFoVTXHqXzYtmG/fTp4Wtrn
HPMgl1KAOABI0j148kuatz//ZvbL8jtnQpdcESUCapfN8KJ8BgpdyBjI0qo47B6Z
EY0eQzGN7xp+pU6PB3q30ukmkgKu1gUR964uMzC05gnYeyJnQpROYJomdtclPDXE
TsqRzrKMyk6ETOz3Jx6d2Tmfx5pR/pwP4uNy5MlyDghCCBHEFAYTVlc3olgst+ve
DKRyPV7BX1/FhqG4mEfQT6Ru/HlUiOKz3dab5voh+bd+e0eaDAYx3tdc3ZPKj5+X
cArY0f3Tm7jMzGXssRfgb2l3T+Qa/djWmmzP7AB6gY0x8hPUZXLhjH59MMah3tNu
QtPM1l9YmU7uDpDyo5NrR3bCQ6mdJj6nVyeYcn7eEGQQPNed54D+eEmWN3Cymvrw
jxRAPKl8WKVhKnNw/B8mnP5bPLuf+tQna8HUTAvnl6vBE/K5Hj9MU4G1EjtgUS+r
RConvyiqqgFsjPuJzdTQSu8QTi5pG14oKt1BQ6L4h0EFbDPDHxxelatuIX5xgpZD
Z3FYsdInEqulsnwd7LdynaS9Wr9RPdxnI8+FplFYGVN6x+OaeQLdMJ5dgn2lZW2M
X1eU8jBsU5HwiCjp7/3uCQX4nMf2sMbQaSbZOBW+e0w0Ww81bVJlMR/i/VwkBQgY
kAftTL3jVkgwWWJfIWttCn1YqgMg0za3XnqvKemeP9ODdvc4pnHXLCDYQXl6VWQt
IFqZ7UAHN46bcllC7M9sYFoieUlHw7eaHEFoNaPSLz4DQAhr6092PM2S00gfTYwi
rJJZD1dGEnvT4DmwY2CHjpNh4VL7wmNcK36PWWzvlDRdmA/8DzYWK5bppeNYbxx1
E30vvHFBDt3qb+IrdWl4tk78Sf4dBTcUB8HlqXCHBK1Ko/htHx7LcJnx3Z/yxG6I
Eb+1lPxZQH+JKb8jzaH8EqBRl8mtyOvSE/ZJC2m1wChjzaUE6i7OogLla8nFcDl4
gVpOhK3RMGBiRYhJFiflZMiYs6bEShTlmM9XsMTBTw22U/m5ZVHHeeDRA+0qQThm
S7m6CgeGeivVWAvRK6xL5zXRXdOcQW0gVz6A48hPZ+aZ7KVnRoFPupGjg21NmJuF
eaH5ArG/F3/TH4+v+rjs0FFrINXqVqqv58disFem7iEJMstUC5OAv1KfmcpsuTC3
Gt7QbrBg9FqIGsu5Ug+ZeY/EFygGkMxUZVgh/+nPSG5wJrdDZg2hscgLDj0x1E2F
mz2NPaXeVd6eOLL2BpBie/d3LjPzXS3Wpk/JdpC3AO+p0pBHLXCTaCJlWQPrb2c5
OBLaMq3KsjD3KdifU5/r/q1pQSIBW25gOqgiXPLHMJkpwNawMvT+TTCDH8hJJV6Q
t6f8P3y+fdHJhNoOA6N0TTZ7ECALB29q7T39T7IWrtMxoUH+kP4N9qwcMr2Q/pdZ
qnQ3q0ThPCtV5Pu0IUWtX7LUuKJp6q3gjLkoHLFd745NlvvQctw8nw2wGQgh6rzI
4fTnZmij+QnNeL5vnQfFiy111uSr3l2DfEb1ETYZQCPi6X89EcdLm7uhe2CKLeCP
WdeT8Nbrph5JD3atMgZ6UocdjaHVAvaGMiYidirZsV8v4lt89ig1dfkTKCxDY8Ns
w7qz7DjW0yF1GXnqN/ipHJGX4Q8vA+sEeSaKTbh17QrCLbXtgIuStRsBv4GU9/QL
qloVsTx1XR7oY6+a+W1YNaFQbUUhDQZ6Y8EkUltcVzbYThDSZfoTr8j/Z5fILbKX
oKUHfPLmo00OCCvkaZA/xaMDQ30VvMSv4FKb9R38nY2RwKGJJjut02gea3qcX9uB
p/sSFFjjHwyOGU8iGYfn4W7cJP9T+xC404GgCkCzBJmz7tCFZyeduCQS3w8mftSK
iJGdqTn7aLXZHtq5soWDWAvKJkq6PO37A+8Zlr1K5zMcx6Zdkp7JFg9pRWhuaxFT
O4NxgleYVF2qunJdHyPwKsohNHRCJNmzueSluh4JomRSdp6XLOIJzINUT9N3lCPs
IBB9WhgECCR5oHAq152syPsysrG0OmgU9LyUAiLtunAD64e466/6+tvAORbhzyow
y3TJnEIj5ZJeMZLKDxjCsBX0tN+Vn4P7XhEM0fjPc+ngK5c5jFbNQDWDBZCzRpDF
5oECUtNWFCvf0Tp02qzdHNtcsuuV8cmjN11+k7Ajsx80EXubyieuGehZBYeQNUwR
+uQ2ZH3G5ni1B+4UZSXi46y87A8RGAtY9GGMqNg6jmzPgEwzE29V0z73i8QAGai3
1/J1VoXuuG6w6a5tFq/VbFB7zJffBmuogk2ADowsZ7nevXMMaDfrukdn3+FloMVk
gGqLJ2kLDK6nsp7lQXYxanOD3toqL252W42WhSZUObrMmy1WlaU6HoEIuRmscOUk
dpjBVXyINC01QEFGFfy5w/dpPkAopVUhvz2C8kkHBpZFmECiXlNs3Hq0rvfwgTwu
yohOsaOdJndunEthw2MPF1ibSppaMf/Kd5ijDOUyNmDZBoB4ImNh3hLIc1GNaLPT
hnbKUqWRaoiC9JMm14L+YZiTMk/rOHv0LIKhZuhG9jaX69bPKFqWGKoBwNJwPVRq
yaGWQ8BSSC5wC77IdtA97aSzBKZJ4iO0VtQZXoEU7FmmXD9K9R4Kd+sH2yYDCVbS
epbkLJqlLGXIoHQGGtkXyyxEL0h/H+D6mfVx/NGNuvPpmtWhKNmqemJbFKaAf8ug
Iqa406DLZu7n+A5+3nYT8GzZdrBGpkjXB9iAyLm43jxSAHqhwXJlhBW1QaJyaGe2
HHiZLtNOQxuW53sCtrny2hpGCelTjkNR7i0ZlGsNR/qvLzwlMEJCFm4XJ334i4eW
FWcSHWaCVEPvy2FTM6Uk9JIIYwCCtmffq9QGwZsEIajMgZm4oQd9wLrFbdtCNey9
tWsXI1zhl0CdJqMZBOeFKn5CquKA+Ues7ik1kAD0yT5GALdNKMIt4CuNnDIPj5dK
1easWLyQCB//JtlZOL/szL7SAgnvWCct7ORepUyPJfyQtmndw65j15x25rhu84nV
yeYN6U5Tpgp2oEjTFMFiy94DvmLfNTBPZpvftS1oy3nruOHMxj411L5ikOn3uMJj
RreGs1h3b0wOiTYQ2qi+cd1Q8xz/l949vrXVU3Ralo8UV2Fd62MKCZRgj1xUUzuh
0svhGuTpkoI6YN9ydQphjBfqwaC5O9+9Lg+g4lq7mR+ExkosDe9mayh+uACvE24V
+8IO2s0JwlqaCOj9AeETb1zWYqATCOvtRnOOi4w695PkwIrnqpOxlHe5/rXXClfJ
OEY8etbxj5GBpDLtmKYLVasslS5eJLj0H/qMLOAZkt5R6cn6k6i+YgTnBH+bRTr+
13YNb0oFpg37pa6V7k5HYmo90L0Nukc6fl2EbPIUQRouO31Ym4Ml24yzkKrVp4DR
x738XYEEWDP2ZqvzNw31f8WxVqRf1wA4SKOmzEC8dORbxINzTxZVWtP+8GfkW2pk
7KssDa8hX05oUh5FDRl0Lzv6RRZIN/cuRHtB8CcAmf1UFvIkwERsgmfQN+w9e4KR
iaGdVii9rSr5eOPuqoThTyRmByqP7I//wva3A+NESQ/fBpqNNheleP4Mu4719ZE1
IyqXeDFcPuOc9Ogp/N9r6z2CEHQDLCo1Ww9PAxsNN64nYZxG5x4aBA8lcgGiBNNm
exBCjfZ3fode9X5d181RXCYmooxD5ETEwPIgd7PSqaBKeQEnnsis4AIEihUqJGpE
PqMFqwYp4Ezl5Ra6n5yT0ygLV2Cv8GJKkdYQhW6JyUursfgY8+iaCBxcPslTrE5b
Xx9cFwKd3mSeqWg+r0MhN8dGZgXqhguCAAHQ7X9OX8oOIi4CaNv6K39zJS/Dlv4m
x0GfNkEIjd+ubaEECYj1mrW1jGm+O/t7IcW6wH6ZOMX+AbVr7jSFEMZz60h8i5vg
C8yBTJLY53zxz8SP9xFbh7JcrRpGbGflIf2cvhD/WIGNPVc9leNAtvFMaEiECUoM
JnW78k3oo7P+XEGr43IeBp83F+4yrBUa3b0JM3lZWcUGv/RjNpMa8btOXIB1+/4P
il1LVyDr2EKPzJYmmCaeHMgSzlDXjQFbviTR39EWA2yfR2kukAX31riHzPjHhSZW
lLtiWT3vpEZrxcs+a2l33nFSYTXYA/froRa9vOufln20MabpY4EBUBW2e8S2v57a
9xkcBVlqTlFWQ4T9ip8UMebTpQBm6x5+ZObC5kF0k7O/mOUVV8o6o2C8JucgfKu3
q2CON5pMEY4qizsFdS79LVEWQYvPftrT9GS7VbTMOHWsU4c0W2lyUQpsE68oEZ85
HYq/hb5ixmrBEGMLgs0B5AnCTswb3D2fB/91e/kzE7JSmOPS42IEODAEHrCQiZ3p
KBKPOlv/T4wgb6EEimyHnAiTZs4olCcaZIFdMzNT99vwui8PgYtmQ4Un0OQRkhjG
YwTsXbSnOFnW+ZVOftm92R0nnu5PfpJ4BwuZeJYX/t+i93HDwT9aab/iB2h4hB9/
YORPs5E4gPMcBDWpTQknKVJ04TZqvvOLiIiLiqmNqR7WKSXXy1BGTIjcSKvmmIbp
qB6ibhmvxLP28ytsq31xblQCuNlULafo39BSmv+A+dS7FqhAOuIEuNBTKKYJNtG1
e46nmhbHKE45VfSRFZyg90vV5LDkYpHHpxFlPPXY3ss2RhguMNPDpqEdr0cWBLPL
U+/TZSzciWeg7uU7ZdZdUnv+2OGlzU6aMLUSb2XC3xPerIrNFd8NPjcFFLazdm46
ejo6WK3JF5blPW+zQMcI/5LuhsFMKfO75wRT28RPF7Nov0DRWY7SLjguxKyiWkGR
GR5lR1/D4hPaGiH1REUk59WSnPP1vfzWQMG2lMX9Y2Po0XUsbUgmTnk5L/MK9j4E
LMlzlur3z2Wuyl9iwrt4FhYTkY/wZLJvVnXfZ2IJaeqHc2Huz8CImyyQnsz1gzzu
5odzNDsMkq7fWZ/eG6zJsaxO+Ylt9teZC0n5QEmYrj9GZkTftc7CHmr8JhSNtPEV
KYHg192uYyeqZi4f4+S45Ll5BWkMaeHaaVZaL9a0PXMwyXp81n/wjw2ik4zlD+Hl
HITSi3CKfhe92/tuk3J1yRVfJfP5wsTO6ryJBTMalpI=
`pragma protect end_protected
