��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�w�����)���F�+��o�}Rc��(�f0��k�A@j�M����=�d:F���tH�|>Ko�-I�Åb"��'�s����j�B����><�����ZeK6��^�s�B�b�R��O�@�� K�)��d̡�ͯ �ml��o&#~��k����}��<��Dz�����>�WRN����gY糖?Z��&7,u�.�cFb��.���� �j��N�%�uM���-i�f����3;�/��*�f�0˸�(����O�yKǜs��^1p�̒'�Jm�Q�w�4V~U �joֳK�m>�#���_Bd;
n��d�5�n����`�x84�d��Nș<��.�����$TD!�[ۊTQ�tC�+n�����TΣ�����p�����G�:��~*�:��	ur�h/[Ri�+��
��Ȋ���K���,2�䓡@���A���6R���\�Ü3��{rh:���ZEu��4���_�J��dz�Ҩ_��N��>?�M�FY���.i�Y��P��p�N?��g�#Z�˂�t���H�����|�;���w�P6���t@�C�h��;8�0\���z��H� ~�P�iy��GuCf���LJ�,����ϜUU�0�ߠ��e�K2u�S������ּ>��H�FV��c�x���r�,}���ϰ�Ӑ��F5l�`��1J.%ݙ|8��I~�~�3}�Ql�g�ۛ�Up�d�CH� ��q�J5�!�p���1=��\�c
Q<�ϛl���@ɵ��z�؄̪��aG��p~�c�N�����rw7�e��i��.�n�x����Y�[@�R���n-��$C��~f���U�Z�<�K(�Ղ*Jk��b���(���
�f�\�_l:x��C|��s���ѿ�t{�x�֬��o�ܮ&�Uۼ�8���#��k�������K]t�b,�U;E��|Yled*��Rg1+LO'(�
��՞�pYR��C�wř�@�#K��c�t�pQz��C".#W�c��"�sQ#�� �̇&�پ�4�b�
.�4(,.{9��h*�q���LO"�p>f�����Z�18�x����!���G��l��G��p���Pyn��A �0�܏P��2���^HҾ�;��Q |Z>�����ޞR gN'iH*W�����I�^�ɢ{*�yu�^��=R��xjѪ�׀����#d{�J;�W���P�7{���6��-�#ܩ�gb'lTrl�r�������8����S¡s"V%p�ڻL��hH˄6���&�rD��f��1o�|��}tDQ���N|�'�_�MTpx�N�H��ח�XR��a���=�i*���cYv�����̅gQ.J���s������^L!gmD���)m�Q����4�WVE���v�G��2�v�TO\�5�!��OEЍ��SD83EZ�&ַJ�P׈��	���g�(��B��@�����w�.B_�s:qp|�-څP����@ĳ���3nr�Ɍs��Q_۲��|�b�O;�z�fn��;j��vq��D��p����lEWw�{"@�䏈X0����'ڨ:���^\��_+k�v2k�F��� ��k�A�kߙR&;��1ҜJ�S^���4��:�*�((�*���@�o�.N=��o�_����	��C`�7�0J�n,S4^� ���!���b�l�HV��������F�a�G��,�!=acHI�Nxќ����� y��QK�t���Ƣ���s�2���^���HoRͳ�&�"p����l�a������6����VNuh	ˉ�&^Lܵ���M(̘�k}x����Al�$k�&վc"�� �Ưa g���S?m]�^��YpZ4��LŊ��t�nCƲb;F"�(�nK�5u�?2&�pT�C�~qmJRS#L����Op�G�O ���N�NR�)��0����,Y���"�L�{3P���vN!���q����X>�����>���0-��L.mC�h�d^������!欍��A�~��
w�������Ή�{v" S1��v6�>&���1��)gX��WM�b�Ey���*�o�!��T�0���-=�T�
? ���n�-��6��A��L-����/�����ӝ����ԁ�:��d�f_�P�o}�̨zu��}(9�i\kAS#���$��Z�®h|�s2B
��
�{�}!Ë��	����cB����`����T*���A�׃f�+�7�
��ߖ��@=�q�@������Lt�Y|@���
?ePe������A���_{�3le�_i�v�a؀ʾDb�+g�;���h|	a6OF�}G�b��S�s�':3aE�飄������Ng�׉aj�Q�	� T�-�-�Ӊ��@�,hvg�ɔ���F���.~;�H���Ϳam�(���Q�9��
�5M��{���F��p�䩷��[靹q�(�Ɋ�'��4mt� x2+y�>�u�ҍB�M��������˨�٤�{���S���C�*I�h$R�=`Ssְgc�6��"�ٸ�_k[ę�K�؅@��-���A�a����Rk�N���j��NP���Γ�J�?�G~���!@������[4;�Zֻ�����JL�аeˋ�L�{��Z�Kx���s�ȋ��T.{����/L@S#2~�@��)Q�}���8��r_Z:&�m���uG�IN��`y�FJɃ�e^�/��j���wV�̳w�����Fc�<�͗W#�"I�ށ�v`�~"DPd:��YS<`�M�[�����Lk�����}�]��y^�{[ܪ^�H��`��J�`��"�`��`�*��ʬ�Q���(����ˍ*���߳?\m4Ĳ�����=��[;g,A^�?��`�Za���e:K1q�
 |%��4`�\s����ۆh�v[T�h_�y*�?�?x����,������ݯ�=�.F�F���Q�:�)�/��B?�����K��mJ�O�,�{�+iW72R��qf 5�zC.p?�G~/݈��l5 ����0�`�WO�myrb��7{�͉N�,M�*�#�i1����8ף����l��VT���D�;F��p�	�`[B+��맆�Ė��ӕ� �a37���z:* �;yS*�~IuH���+���1�->X&�wΥ� �߯+p><�vOJQ/HaU�	�����]T��k�q����	�M�3�.��cA�!zLb~�R��<,j0���+	�90y�pjH�5�B)����˶�^�����_�e�\�����V��S74�V����X"�o	�[k{�A�>�|���h�;uc�M���qIh�J�Rwi��f{|Yӡn�e�ǈ��	��=��o�@�:�H.@��4 �9���ns\^	Ή�]�n@k��A�am%P�E6Xf��q�֜nC�,&�e�=Ҍo�����[��i��d�g�~�v��5I��7���Y��"�o��Cx�b��~�1�+��7�q��N<\�ʣrS ��Z��VY��bE4n�ߔ��7�g�q��f.���X.�5sg��_��4�sJq��5��Ⱦ$�$��G���a�"�b�	
:�!�x3j��u6�\���P��\ ���}X�� G�k��c�l�l\�) o��;��[����O%��@�irVI>C��y�,���:Ϊ�S��}�ćJ��Y�B���-p��Z���h�z���O�]Ա��f�r��f�j~+!�+���ۯ�$�WJ ^���q�\�f�H6����)�{+�3�D��{��?���<�^�>�5��\��j�BpG�}'i0Ɇ"i�"�A��hg�|�~�s @���&
2�i�Ha꼹L����7��7}k�ɡ�.��v8��h�"C�.=Go!<�f��,��nS�.��0Ψ��$t�%ª��fZc�"M� ٕ�5P�'eL"}��L"$�^H�;��$��T}�nNM�w:��`�F5/;k�v�)!_���l����x��ı��_�#�%��vOU1�&�����9�*����-^C��H�Ԓ��[�-���ck�]��QNw1m��o�6{Z��%�`��0��tw�,M�g�j�7Raq��O�$�ŕ�,��'��7�3`XSe���b\ ��1��C@�0x��/T�1����	�[�\��eå��P'Z�G�@�:K� �&D�ʜ���]��!jr�6��v�.�X�,ś�ë��rȉ+0d-J