��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m��P��R�%�A�Tf�/�`|h����_���c�h���<�.�9Dǯ�>����{niB_ڍ�"iMC����8RP]41Ǽ}y�!E�U�+L��O��q\�Z�O7(�D���3�!v�1Id��A�a5y���@����k�5Y��lIK��vk%��S��as5�Td�?t��Z<��OڔX��`U���\�ɶ~��~���{�����۰l��d�2m�
�`��U�y�@�M�QJ���� Cl�#g��u�$�W�< i1/�a[}Gs��5��8W5|�P�)kK���y4�}-n	I=��A��K4��mZ5�!|�s����oҸ9���m�iSxb�O��ĉ�~U��A����i/p��|2��b�wWDP?��|��m���(���\�Ro6���˲6�CatGXe}��b��"������������6)�z��<�V6�$Z�J���#�X�Rٜ�F�����{����	�B�q���L.kE����j�kb�!���P�*��:X�	$�.B�.)E��
�3-E'����i��-�˩��rN�,�o�r��ơj�8_&"�i��h��b�e�l84���2��kd,�|����e�9�cc��R�jv��@�zoP�chR=�4{�:"4i��òY�go��.A�=ٽ���>�4��bjz[��)y9x�,��%NQS��s�ٖ�� �x$���¶��7_���S�h�}̈J�Ť��w��bF f����U�EE��������J�*��yJ
`�Ҏ��;�N�H�*FW�ԕ��ijSM��ڏ�\�7��W8�	��#p��I�s�2�ǰ�X9�b�&P���AhԶ�����U��1���|,7��$W�e�1k{�w��y�ʁ���TM�ɟ���]G-տ"5h����c)�F.s/3PbE�l��d� �g2�����P�B��ȬXZ���eVsB|�������J<%w�
���ǘ��!dUX�Q�R�C��E��[z�J�����>>����eą��(���Mn�f	J����5t��� �̯꾕�n���;
����B��E��O��6�c�V���<G*��?�������\�!qj�A�&P���!��o3�A�EEC4��P�IZъ� �h��J��BָI��#�zJ���c�����S��8�[��l�0�e�a{���HX|RS�w��o8I�Z#՗����)n�M�����j%��؜N�eC8<�����*1rr���l���Z��Ig���>>�I/�� $�������:��X����o8q]^� �7'���1d�s.�@/|����[�ԯYA\5g^�i"ڸ
Ķ0��g�ǔ���}�e��1}btf��vZ`D���Jcbq0�q�'30��ӟǠDr�?r��*����daM~���|��!$����A�71��W���C�ʃc(n�(���U�u��|�Tv�^S��q}��t��ZP=𿺡i)6%P�u�NN��&$ʰ���.vV�c���&@H.�LP��Ɲ\�p����X���J=���;i�e�\�W������K��}׳�R`>���_��D��30;�J�
P��rI\C��A�.�,($��&��Qݙ�]Mg�7qAT-����̘��1ٚA�� ��~	��"R�*����;��*cS�T���kl�<	���������]���~1 ���t�Qy��ԐQ��.\��N�/AO��b?<S�a����y�BH�q���L��_�Uڙ���sW�bi��f�!^(80�'��a��莑u"���˸�?���%V���/W>��E���#����:VG��Y�M0]zm�Ӥ\�s�݀�`�I�G��?iu���)��u���C
���IK��>~�j��7g�F� *�Od�#������
@I�1K�uX�0��f���Xw)����q�r��0clDO�KQ�6K�7Rp�?�9�m�n��ev%�y3���d�<��w�c�8)R�E�onS-�R�u�����F�|�ĺ�}K��+@#��&�ߛ[[=T�4R�"��µ����Wvr.Ҫ'���[�uI�.����/Y&�	�cx�U��A�Y��Z̙��KM��+a���<��a�<�dr+}��6x),�G��C�]o	�}��ZJ�e�ꥶd>����uJ_k�!���_%���:ڿ݋�F��-'�;��+�l���pH����S�.Kx;7K�9��)�Ы�V��LUz{���5�^��"�URT�$aE�'���1���6(Q��E�?܉���K�����&{=5�&w�`�s�%Baz{� �d�!xZ�'cT{�)��/ ���#��Xы�峛�< �ьj�	r�a��8V��``�O�D��B��]�D��Pl%�7��PT�?ޓ�y(��.>.m�l�Y�X�+j12�@ {��@�1(�[�N��y1�&���i=u��3&} �v�O�C��	����7~z���i�QO��&#�(��w��Ģ���'�I|ʧ�_��j�R0o�G\��t��kp�WQc0�9s����w��MJ��HR��=�iB�Թ�j�`{xG�t���ߋ.5+���TLSQ0��o�"i�-R�R��<��C4=;�V�ã:"�HU��"}$錿����-�ΟC����hcɁ(��,u�w	�!(q�F��$�l�A̓[��սiD��a�����(B�[��4�C�&�J���ڍ	��x^�ܚ�+F�f_�t,����:��ü�!�fo�� ����Q�K#�����g���9��*m,�6E�<��"�=��I�і^�7pt�7Y2�D�	]��"��(����[�1$I��(�I�d���IfHﲎkpHM�G>���}���wu@9q��`�Yd�W��������?l	΁�p��*��ؒ<v������	�*���M3(�~^�*����E��� k�`ux��Dt�u�?�eU1Z���"ꓝ\3����xf��}c��v����1�GW����h��xx��+M��9���}�#O��0�KN�l
����MuH��t#����52'���*�ͳ俿��y9 ���4>3�hx��gK��5akn�����qb刵�a�[,oB)7�F)�!��;�.!"b�3|�������X'�m�� ��zG�|?�mi;�b���=��&C9�^�U�g���<�֕��{��OT�qG��S?_A��s�X����G�QtT��'�<9E���+�ܭ$|r��ٕIv�4s*?�%&Q���������QN�ѐ��$UB�׍�;��V]���m|��%E��v�}�iW���g���GXN4JV��{�sg��TB�	��rK��=��炔�9�b1>�u��F��sl��8��I�P����ތ����7ȖvDm�Q���wY%��W^

MxtЙ��a�D���l	�W�hKz��&���MU�/3��R�:�1�R.":"tQc�nOt���V�`T9n���O�OW	���[;�!%���Bf_�"��\B�);��3aL�5�$�0Xe�B5�f�ȟѳ:u��M��xml�%���!��h�����S Y�x_Q{��kq��2�/+��RNZm�<�x�]2i�6��=�_r �Z���ym����!F��02H.t�_-0 ?(l��N��j7�s���@��W��23�����OQ;��o�T���^��%��NMho�T�%6�*�\�$��a�^��_����:�c�Ō�p��H1w�'?�wc��Ӊ�Ү!�a��"H��]9u�sf�L�����fz�w����[*��iN,�7!�4zkc��NI¯���Q��I@�Phz�鮒8-��cE�pNHo�)�f��9��pQ�aźu�i=l*�hS�2�2��$yG;8~�{{�/�J����f
Ln�NҫN�so�L�{���Ъ2{��:Nd��)�5%�(8#ԗ��DW�9�p����eH����H"�8R�f(��/�7m~{|�6c*��صҥ�I �/(����Q�C��h`_�έ���D�u�<Y������ґZ4�� ��hFt��]1-�Z���4�Dn�+�N�z}j�����?����Ar�9���v��6�Ƞ�oQ��%?�n����������~����3]����z˫'��ݕ��|SY��Y�D=�<M��#^"���m�&Hf��[s;i�U����2��gKpi�|��"�A�y�~����d�