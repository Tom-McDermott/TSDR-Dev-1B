// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
33I/JuUQgItBeAsiYWTxhAEbmkNlgHORgQUyEWJEH43nPzzc3MLqIRPgApBzkicA
ydapXpFsiR6vltZziUjta7OG2LThoiuCF72kMr8KQdiKQDTu1uGCVL5lBr1Yu+/i
PXFWLYrVa7GlsgJzb/pCem10aClSunN3fN3Udu/5bI0fGTMYQvRdag==
//pragma protect end_key_block
//pragma protect digest_block
mXpbu1zCmgXlFyEUk2MrAcmchjY=
//pragma protect end_digest_block
//pragma protect data_block
fVXhZ/EptOeUkm4DseFk/TDA3PgHc1g2wr7ipjNRCaMZA06lEp188hdAwCftt3+R
PQhbOTAv35yPuJpJvdJchntsdKPlqSVi8fBSGEuWeDCJelFGbbNyE3cVN+BLwkiv
+1rxaZdqTKC+v+AYcV0goNOpC7q7FcV0IawXdp4zh7oTSSVIGYPU9lGOdIN5gl/1
zYjpGtDXD8+mhkJKXPseKfJaE1mUiLF+kB0Z+SA918UV9VWJY3Mq8IzEFTijro3I
chFAWSmrLcp72GUKC/XtmpVNqDr0MhlLB1utm8x5BTg7T1/2cZjS1hVYiU5z62mT
jQh6Q2JPqKaKNJcQUla+z9JNhHFj7PQDAIZa0z9z0Pb2ahE4+vutoNAQ7thUgvv6
UXpesE7Ci1T7snpRhxWykRU7v7cPZeocx2D3znx0TpNkbEuE9rb5FoE7deLstBnf
/AeGwhpgDuWf1HgqcspHlmQXwBrML2u9+QcArElaXl87p2tavPs6kWDXb0DSSzR0
4OjFGPXVktFhg/TA38k0iaySfROGcY0c3/1eO+LdqGwaE173zDlvyEqGQsYiOoH8
R/cDlwk8XX8dH0Ac7y+CuLdlIXr7zm2Q/xxW4M2cnQELBsPGEFCiXm9i4HnXOsS5
RK2rU/REFxXUChAUQ4XiRhbpAcmU1IYe/8vpKh9xLVK/mMGKfC0/EaNAPzYSjCmd
uLnFGpbDcgWgaawemLSIyACIF9yYdc31fIwobhi/mvFH8GfDuV2OICybUIW8eYqy
2PBiqUMYPuJg0pSFGdM1U0Uxv77qzxzIspW4Z2ane0NuOwV7L/2yvnKmCXDzX2uu
3AGXd4SzuHsvspWhq5d3nvXGnqyJnCQ8RTsLcniJaiUS7jz3R13CNHL4759rvU/S
Akp5QbcUCI9VlKfziGYY6ic5f1du8yJ6kBvCRrJPJ8P5dgWrqfwtbCc8kM+N++t7
Bvfi4km/n7wOKRVpWJ3DagGzUTcp3tNUwhlMzsMDd5RWTCXfHNc6o3dmV+CujoX8
r/MRPBFdU1t5iiQ5oeEbzvrmRqXV8hxMiMSRsoyxp++bWR4alqIgNaomliecqEiZ
NTg3Mx9nsGOd2zqN8h0JlcaVJ43dk+Zp5bwqeqLv+OvxdICl7lsB1U75caFcQDBp
vFjMq07fY6d8W71zwG4elDb9JpdxlNxGhmIFNNkmqsQKkK6lEv/wsYGwm9vu6sWJ
1/+r94Wc11pVrk3jG3M39HB6aPwoR8lAFpbKj/cet9gCWTPFmP8Kt64i9UAHPsg1
k6DIzYQtxK6gJHcP7IsNAS3oFm3NvGoVVN08KKGfL0HVwaO4d7f8rnZywRjcpqAN
nkJtolI/NY4pT2L6Dp2GWYSeKtPJroJMcYaqvKPK+nOxwzq/0gDoS7FzlH1F1LYP
m1YMaevQNY0EjIIpM1gqvJ2J3G9v0LWox+3oHLYTCfInkrD2mzJmhDjgdSn/OQli
wgG6v8j5Er2YQuAcx5QdxG6V/TbQQ2BOjBUbFI0sVKkuZ72Eax4H6O7+XOvVyV9E
sUn0EOwKQjevwCLkMuM9I/yHjhsBWjsHmGcFpz0gBIq9yaQUkpWMNX9pa/yf73cD
03E5iIWb6aP+rCFej0fuOj7blvg9ubele53prHCPPERRau50Qo678nG4yKgZXj8G
B0b0wZlBtVoJoDVsyf3d03BTQW7duIX4sZiZJl62bx6Nvp5mxUeob3koRsOJwUc4
98rbCHNgs3dyz523u+Zu2Wcq2X443NNHbTlCErpGBZ6MrUd5ySSoToVZT84SRE+I
NEcLnse+LTMoX8K45s8+Je84iSTsj3dGeB2GFxBwGA/RQVScBNJpuTyP5Kh2ovKW
JM9BnQc5BS9ekdbZ7YCpnJhN8aTMSizBq+2wPITYSM7fazwb9blaeVwLTxNsGDm/
s4ZlW+OxnOPzzKtiaXhuz8zdHKqMMi0FyDtiNhrrtMNmKI19cc6qTiUN3gKSFVCc
tXT/tHV3y4x3xWktTXo6j6ebdTOdSdwKpLkX5EwKJTjlZj42Y60SH3pN3YXI3tED
cdoDgQZEUCQcYXjHKdnFPwvPNJvjodlmgB83E1HPs7Usu+AFtHDFFxScrsAtBTSb
2gHSziTBSw42Qc4j0sOaMi7u8OgXUlqDU7yUh2pzpvIIwahvBsdpbxxDZ9JNhh/P
SvjtH+Z7JcfuoAEM2igHSlSxHPqL1UcCod4HBaYggqigXlBC4K0t7SQB9HDM9utG
JxS0/D+bbky1BaP9xdvymiGOHnkx7AsKm1cNCcTfvHEGKvdQAwBllaRREKWlZLd1
U2loubs2VT1SmrL7/1CamTeK5v4ppfDCWnYJJ58+eSQXz2GAnUuyTz7XLEajFsPh
meeYYlbU8ub3f+bKX0rXHVz09vy/jZ+WPa+F7fttRpnNj/4wa2NHvdG1bC/6qKSg
SEbjphqzMXSMBBsFXualApYlXY+uzfwWPJvukh238hWGjDettNaUVrBWGTNCjeL0
7KN+Cs5Bquh8yXi2g3ZtahfOPitC/vbUEHBihCbn4EAcVNUreRNE7tON14PNQlmT
/1xmHypMn11S1yaWc/SsfyUpoq1q64J/tW4oca+vu2LZ+U9h7c5dAs70XxudUAHs
JVAgxXDaP8Mn1EALBk2nHzeF2rUqRnVJEW0XaW8mWeSUg8wl125rH5ZWoFDRiKpJ
hrv8NT4W4X82tZ4FR6SLUKedBsOOUicDg/+tqsp5wSo32FuaX2b5IHTKnj9ovkQA
4pPilL7KzetHNzEy/PWhjio4P8mDky1QnpL4UbyZ9htWx2QBV7PHkR40Ci1W1kJv
tDfyaG+7vzQOJAkWs+Xa7ssfdEnoOmNRvdGWU/NQ2oHW568SgUwFDN0KHil+QNXz
r9zxye6j6u2nGQAuoQI3rwCzA2UezpXQTAuiaqAppCTGWRC6O1jVKrXzkDSk/An4
I3FfCr614V+daJ5LULX0czsGjSSqmgHxBhT+vErTYH5iXfizOZEG6H+U0esKHx6d
BZYEHn+SzQdM46UcNknvVSOu5XAc1qugoBWJimEqSqpA612XJYBrmsElySguQDt0
YY2mqkhYFlphHfAX12MnPOkdWtutvmMva6fs5OvzFX+TClBtPihpyzm4GjwOTruo
CoR8Xtph0f6ocTkRDlw9qfJgyvImXGiQ/63Sa3Hv+PSJ7cyuzCDx9G8LQClWw9wo
cS758k50vJtndS5xFtwXpu/QESJPC8W6RYA6MJJoqA5cMnKWY5CXf71j6xR/QaUI
tSQSLr9ypaKMe/CcAYz4otRa0ZXjGH2oS2xPezz/YcbzeKfZsjdShIHQ2DzmZ6gN
8U+OWvsTLZFtRCPTgbNzTlZwW2I55b+NcO4UI9oIOx9EGv+TyvBDFDQTsuWpNPNC
DYRfcJwBviLKHfIH4lBSImMnnruyXkSfSC2R/ooXvngTjUmhfhF+p91+1IXhp1gd
pkPpZEsUUiesYnoD1V7ntt+YRFFKHYtyXBaVhgszYIdFb4YDi0dnAa6w2MkRu7Hk
0E+7GnPgVg1dFWAsPySdd9TOxw3y19+YizwSUr8WfwtJQqp+/AVjWU2Ltes9V5Uc
oN5mD8DXe1lpJ6Yfls+TIAYf4L49QGAhhxQdQQJiHS7qwRF3Ug8ZypAZIKd56naa
Fcr6zdJWi05/3Zd1hEyF34qgvww3lu6NPXPNp7svUQYwF9RKQp48jMLUwDfSejgs
xrUmxUIVnd+DBr5If3wA8JVZSag+nbgKAAqP2Lyi0SUtN51+Fm3DsgzYB3bujfOC
JFyCLFEG1AAJnKTCpMja6YVM/Oi8Bp0Of2g/tseNKXB5nEJnKaSAwgNvS4FqAwfR
6na3vMnviTs32pKp+s1CVtaMZzmxEYHB3pEjzmWlgsRDMaUR8x6lnOFb6uHCsZAz
9oOrzpksC7qv+IfDUSn3+Y7vf92ZFtFwyMZ4gg/qnEANsbGzQMuqOhQ+QbF8mGWn
3BcjAKDuPQvQ/MkrjqdTTsF7f3LoWhFGatSGxvkA1dDHCK7vJiN+tsmkSr5WrEhl
HHNVegmiFiLaxoN2FAfvRJLdgppukQXSSFKtiHTusHjaAptDWFfARSkM7ozq2Jy/
zw8argnH7yxzmaeC8rjLI5lBR5LkC87PsDCKBFTTkp9nRGJyVGriqmymrbc5gUcZ
sZ6NIw5v4xGD0ahh3NPMB4YMu7VoYm4+yZdawdJC+dRmULLZNqdqe3Kx0XjqMZ9D
sjhLB3CfEW2IS32CC31RVof8PyD6TbtW8pqfYMSLY0svbPlKdUaO14EC+lWwBNus
HreTHm9EJxEyWMYDIS8TZZsIpo/Rx+e3kdG21jKRKSHoNDagbxcqm+dLP2R/pq5d
UUD1lfiO44/4/UtyG65My8XYuH+NMX/FpAO6wIE+i0Wgj9pEI2TYF60w2AMuMHwH
qYDnKOiZ/fxdejSZWt6ec0TWx7f4akaB71S+6sC5wGpZ/0P6EGc8CL7MuJKw0XWc
sZ0Df82vATW6OQKuDcTdhGM5C9R5VeA2lhSIXZd0SnvTU6BHiB1iLgK6yHyCiF+F
eD7XNGdVB0bKO1vzlxo3ErzLX4YUilhJlsiMksE71AgHbwmmVPfpPFyqnmV1/NL3
ti21T7B9H3W7Kc0EwnbqkTko8aMGordUavjyxE2x8C8ZklJXybL7rcF9sLJ1wv61
HCJiKwnl6pZDPtb+unXw6harYzErPzyUPTPmo81zXZ5+zrgXMG3JpTfdaqTJ3U9c
ZGLLYidWuXoV/TUV7EvBFpkWxmRmNXRjA3DAtf2liZ13pbMsp1XXRLFXwuRrGE/w
1aO/l8rokhxAAR0RX12DyhVzxTEUK1Nnw9Z5lxrMzoVvrkbY1/IdeWst2wm0CdZo
+GdjCO/CoDHcY5HnonvuGL7YaM1oQfN0jC0Y737D+QqHfg031YD3josLiczSGuBt
Qe4toN1v42gXlJVN8ozdyCWmfH2WdV2L1Ewp6k1Rslxjt58DwchYJnb6RJ/FsPPi
JN9jxQDnuusc1acN/FBk+bFajSqzkMTziaSCZKjFm+U7dgQqsy89EhLBuBd9nrJK
CTlfJE+5kwk5tBWOs89LbjymoWxjvagDwxSOpka/Tr/vX8gR6ZM4YjjrnBnJEW8O
S9a/IEnerMUcd3BedI2/eM7FP8ye9kj5T0FKEtKb0Vcoaoktf8o42nbYoJ1tgbY1
JfYct5tS10+U4dVzmTIlNMpIhAOyJwenzAWdsJiSZeF7QCfY8Pg330Jrh2N5ml9t
FlS8dDf9+CU5EUg49T8UWotJutgPiDBCDXNKDRu2dtLNZEtCpUlN13Apt2dmrZjh
M3uABOh31qQjdHf8eP/8cO+4cwuVVGpwMVCKAcmx60o2G9czmmHEKS1H7hgVj/Zp
PvxaV37rKq1qgf+eRKN2Xz/yFfYCFdZR+6HWmopQ82L5skHpdOo5tgydFVMqBAwh
QfrB9Lr0QDbAudxMEmPLxHR7MHrNnfq0kyZqyRkuH1Aa+OGkHYMdghNn8JqC9xOE
U9Zoe1SGOtouDLe1gEgr2hByPBc5G8WhseqmLdMsIWhJAJdUnRZbQZ4lHsXvDv2k
2F8sYgvyIdw+uHnLBASlqBWsLjXS3JHnzPvPBLJiLyji4ntihDn8czTC/oL4qGqx
rDrEkv1Qz8ND1XG0mbvBl5yZZ/TPn3yYTWin8lfpX8fkzSK+x9TIgr0jkcHJtf+y
2MS+IH27IzMJrXfsBGbgI2dXvRBwznTWF4kUu4ZqUB64IADrMZN7j16slhqiSGdD
tVWWXWmfvjp3ei337BVdD6cVHjhIA/fptoRowxDxdqJM/E0/zJ4TQ9vZsPczv0Th
Fvqap/iWgZovmLI4UrBWnCYKVGxT1mbBgC9TgIE10KOhdXNCaPsCm7y2TluJdGwU
IezU3KSrGsOCjGSei0lGQ75RKtebFkvPlWnSV6mmcaCrXUDv9SeAA9F500Y0C/ed
vLupJXmhShYGd9O4WPvgQRQXQTRIFQzA/6MwbzwfvHbS+ClcoG376g+iDBOSjCKi
6doVJZ2YxjHnGEEZKp3aqGLyg+RDq7Fm0EjiRysKQffnVwInvOUy78duP36dB66O
cDVsc92shm6qYb3AaHeeBGprElGOKugII0xnKO/5GtiVduaYne/vsNRI4ZxYStWI
n9Sh6ZR4wRuah+3BX5ujawNgf8G0r6U0lezuU/TlLka816psQmPM7gzWhtdEdqgN
Bh2KgxHbcdy6e/wGpQcwWLImcs9aDrMUoVKxV0JqCACR0Oj4M8hs5l6VZG4FCa8t
GB9e9j2hwocPM5FFYGQY5jJYgioYv4mGxQttK98N3TvMJmOMtkiaQtPZaT0hxqGG
+id29JEtMzpKK2SA4v+b25YzWQ0EwPg4IFZXum0B1hUzNlF273bgYtLrZbVWd8Ai
ZIK4z2PztD6W+8XM52K5fEOqEOk2ueOf6nKGBdhsKKF9W1NNmAgzzJAZ/Wo1hclF
DJR9CiNs6/6Cv0j+aFByXctgHtlhO49ztwXa7FJJjl33JHW7Cxd/sGymoEUNnLFK
4Scbno834JHCM61aMoBpZf8gMBH9sn5/jmA29XqFhxrJAo1W0aGtKClBcJzLtzJl
nu/QYll9KOS2qKCPE/qARybpl0rjeVSHHJC3cm9X5/Ah25DsetwzNZ0XztBPLjwB
45sQptH8GY0GydhkkUgC2qECtfFKWSP/Z183fMyORgWKG/XCjAXLeysv+ZZnvTqe
V3AbHig36E4NF7VQZHjXzQ5PzDGPi0rMysnScKhiJM8HWpKc505WH8hMHWA5KT+f
p764JeLWzh1iL/SNfxPrrDjKlzqOrFHFjxzWbWTIPPKkMn/y0VKZe/MfBvIbH1rT
EVGu4ykKQgaqYtkVNN0uUnNqG1Mhc6DHB6GHT6OZpHqVtz+w7NARu+HeenGmxzn1
h5FftKpO09C3H52xKWrhXM10xWLtGiMafd+EJ1WF7c2nEL8L+3VwK3FkMFaYA8XT
en97Y0VPT1fpR4SoiwYolBCN068VYq9LG+RZWRo9r9mYOaGEzSymyk3uriw61oke
Afsa2iRxPPKZSEwUeFuiVGYHBKycDvQN1C4QHaO7U7xKyKSJWUcGAdK1YG3Yb/lZ

//pragma protect end_data_block
//pragma protect digest_block
a3vAPkZzzs88V3WOdVf//t1geQw=
//pragma protect end_digest_block
//pragma protect end_protected
