// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
FOMuKEWW9ctPBtLe09pKSeax5RcnH5QlnRC3ulZYUvNCyIa+kCdeiZ7NTggGl4Lt
GtkacgnTX/BI8oII70WfirmHeJg61uLXfr4YtBhKhQO+j77p+R1gPhIYq0SnoDMW
lnjZ8+pRZVrjQivHKLRtwcyk6HJ6q2U/Gn/s0Wt7B/PUWOqRyHeVfA==
//pragma protect end_key_block
//pragma protect digest_block
HYdTOFJcEwUf4YTLaDn/RXFyQLE=
//pragma protect end_digest_block
//pragma protect data_block
0kx5pHFbCBuGYxxYA7TgCZ3l9mT1xf/tgDugopJ6BXQksHGcYgoS8ADrosZ0mDVJ
Y3Xz3us6M0MyDlt4+TTe2iPcLhtpVee9NxBjh+S3eme132IcfVsqnn89VYpktZCv
QZPcy9o9CmDWPIO5SbOp2mJIlJlnuzSn+ZJQUd6eg1wq7qmN0AIzbccGlrMp6Xvw
pFXXABMRwFQTx+3GHukqhfxpqHyR/XwdsTiOAw63qT8Z9nxbkvYu3+ZiK3Z/q5aK
n7S8e+waq79gRRFlAw4eC6/pu9M077y9RwkjRFh7ClkEKcixloMgOCTRNU+po2UG
sx9arHNTrGxSohBpZ83KZHdWs0NCfqwSz8m8MX/RCFqt44x3Mwv956oFOfGXffRd
G/T82RLm5eCvHw1zCfFJeIacIihwPkFil1NNbqcXgvYZBMaGM9ZcXkrBqtUCJeCZ
pkd1jZG2tyRRa/gPM8TPd3dM6T2iVEhbfpcoe48dbOIYnifw0jNGV8wbmP+61sh/
hA3rw9EwRoOLC/HqW42ZjgmogXrYBFj8nrNw5OlVV9rPcZwv76J0LAdu9JkTA9e/
sqE4HC+8iIehdFNNuyOpik+fQr33hEyBdoCogJBhKEVoqC+/wRrtShq+Yt7LkvxB
RL0XkyBiiYsS6q3/GQxCTa+yR3SHj6lVHsNyfoi9p7sYkBFShy/sqzycRA0Xs2i5
/oTZHiVZpnm7ULUnjeArMEW4Xpk85Q+/lh9sARq+gYZH/C9vrl3sFjt7SOfCi5Za
cxX7zrSs1g5eW9HjIFq6z+xEt/OcfDHq2eZRjiE0JXF7XyKIdNg8dyqTL95eSqOZ
Br2ipMzlZa7hhCHn8tyPPqjm0iWfJsu7sVhqrWwZdVVuUL0wwrXNui9U74rLjkt/
zHPasAusLD458Ra8kOjpzDy/JLPu58WgOfrQw5p4mVNzXnUpUQH00v06EWEhdRw8
vlO1ow74+PNgLMyMtR4PEwQVu7TRyfz4vcUMk9vfmOsdc0a3io87qEEx9s9MFcQI
JnCdhfwB1Ea6nPqxpszUH+VXBFkxnU7ai8nlTZEeLR8CkHwiyLvTfwTKEvLrM6TB
wavF+agYK5NylfB6TjC7eK99RVM5x3FWQnlEQFhIujXFyFjwBCDhQFfRVdmydi3c
vAIVQJb2WAEirYekSHn0QOyNK2rxpRDbrQIQKhuFGgqq4i2iEUH12U65iSGzhUwF
Sddx/bX4rXiH6FTbmtbWhHcfFCw7AyGuB2x6NPNZERcuy0bnduvPbVgsr46H/z4j
EN0WM0FfroeYq6e+fC6trU9h0/KZ2U2jWROdpZBCXZ9ln/d1tvpA5eXcs4uyhA/7
9xjXTdkbWWH89INi6DXhfvE2ZmDcRcnOLC/V8OhXGKKAHfafjK2dPTEUWyVP04nq
v0xEPiBuJJOOQo8gBDNT0AA/yFroBvLPQWzjQEGNGNFb74eCkcMwJPdQ6qUk5D9H
0Z1fD7AG4gi+jp6hC8Oh5nGUz0hPqJfOBE/HGsZBEfWoNGFW8Kx8hTb1GtEzPOq2
jTUQjNspnLGulOifL+NEy6X21v/9EFcp0Lb9zp5qaUFb4BLyoUF+PQV0vv71TVFo
ln95Av75XlRJVfRJB/l0viJyRZ+aoNAdNuGI6GCzL2dOyu0JlO599kk13L7hXPJI
YTc75/X3R4mlD+vudyv2ZFzLmCz4t5519IPoVJRh7vbQENtKxY+7QlKBs06DOoWr
EJFqvOPqhMQfftvXcf/wKda/9zPvSxgpriFIMjYWB+J748aIKcJAL2XSsX7/LLof
zKOaCs4rCehLX6QbMdZFVkpIWJ7ouU+lx/xfVGyON77QfD6VtlLnWB6HwNjreIU1
cx44qk2QljHuo+Hh9DkcbvMM+NgSqYiBYR3JJ3SsIXihjgJlzWSRGz1pky5NyO13
OOHbM3VU2Y/Cd9DmDZaXkdnAyp4wCUzDcTC6cZstDPr1s+Z9x2SVvmf0dEiPfxNA
an6r09vbpT97rVAUCoJ+GDqV3uavv8EhCc43bgMVPi0ROqFWxYr5zgWGVEhMNiTx
tq79AP6vbPDvA3dQbTamhSloUL/Vg+UiPz2x+FZMCrpono6rFkNPHv/KApuNJYKb
i80xADUUaJgqkY2WkW/vlnLhCvL4+AKmzYvjfvgfVs+avUdjhNxomuGbIxh8w6Q+
JuEEFEGaFyO3AS/WpzBoCyUKWl+WYah041JY9KL+nPzCkS8BMslsz8u9YUzHdRKJ
g2YOkLpLN4p1vpc/PsGyVWmoV8qnNH4dBJTz1pJG7I/oKahSZF1bOstk8+F7b3mo
nJx+JiLeqEeOtqmJ9v4Hdt+1OWlBY+ItpQzuT6AWPdpw8jzNU6UjVXvU29NJHMcQ
J66UdF1QhNMfRT5E2kfDEyZun2uj4i5CiVffvvL4PtoT0yMNA2HGgjRwt0eD+puf
1rMWWKa6rUtHd9z7RTH4np4zA1F3ZNaS4YrdJzRi5eYxKOzW0P3guERjkWH88Ot0
XOm3x7mgM0uPFH6bOVQajO1M94MhitCbRMpmZusfzOM67qVCs06u9A6XhRycgld+
8MUwGyy29Q1u36yBJhHKekbq/UNSCZBZBFHli0v6EW6UpWi4WdLjZlIgh7ztmyxg
gVRMrLLwKhAOSNtJkOorKGQlAx4umXAnWrMKTu8TzZYCv+BLYAGIWecRkUZoX79t
oZhG0N5IsIouGMBzvkLXHLMNYsr1B5Zc++psxigIxAyulWkIVlsoOyDemGcnyNLz
XbbckleSCM1Rywz9vKZ6/UHTTeU01hqBCU24G9eFUu1doSqfOC+EgPcDwR3Lq0yJ
mXkPDjI7sTy7UvXyI+zBPyHv4P0I3u6HUezimY/jnh1gpVBL+PON/kpQlTqM6CzF
qiwDRknVOLxqqn7pLvrl3MbOu2wTczGl15bDQjsSxP1CAxm7rMHoqUxhyw3xB577
pag90KFYBHJkB+pniJOrE4ubwiQXsBWxWVQl/nYIy8MN9RxKk1b2NkNDOYrZUEYH
uul2iehlNK0AEa1AooHh+axrsv9O2P8Xs9jNw6NznxQ8qQcwAXIpiLUdtcx2+r8I
6i5+R0/uAiQ7G02A7myW8gXgkslESkAG4/Rh3VFjAhiJQBYNq7ThBxtPw4mmAmJ7
BEqrj2MDbtBg6e9ZkJsawxoCRjU7UmCtYcr/ifQs4fd4TFcE0F5g6F86f1De43BP
247U1oiAryuZNedhhgNkG+S6KSaBfJkbn//pApU6Bg7b7dCHhQ84X0T9DRPpP9u5
GIomaA358VgSelHnDAQzyI3rCDEAsSrQE9UUe1wx7fh9mOhCmrAIIJezxSSJj9EC
Df0K0lwSbtV5uDCEU3hp6vvyzzilUf0Q1doZowWSAKfBmdjKSaNbKJMl7nUF7VaW
bR6nhM762czZ5HQ7e1+a3PNKD1ckDF4l7USGCQROcE9mdQWycqRhzzc21MMh76U3
NAgNUDQ9hPWVHCb1Ohcft2xuxZWlKHS02CAhLGJGqDNqXvBZB89SQE7ipBhnAfYi
VfrroC6pe5cgYWBHGvL84LNGhKD8LiRz5zRdE3xGG9LiUTjXiiuRmtSRNB9n5CWY
xNS3Te2fPaHmqBWMGknpB0fJ+nnbXnhI9+HZva5/Z6/fBMN6IUFF3kFsfNO8PEMc
LxEys7iutTjdP9NWHmFs9rC1d7aln5PQo7i7/wmZWLspgQKOHFapL7+N7MYkcLPa
0sToOgQHAnGjeSE3i31Kg82dvHFPk+/52tI/54hy5lUs0RwSWD+6BWUB+Ar3aBOy
2MtIZO1q1S0sN9g0ZwnUhuriDUBshj89oIYTZV4N1C1Il4njRFazQAvoLwmR0H+m
P+jbhxxnL1D2lKZg0g5n7F8UagxS/JMyDRhJZ5LNg4DcoQPwAgW5o1WIy0HCKFsq
nCpF2+NGy5fnWS73GbIDFwmria1MrCZX2Zy3kqBJIfEHwgr0zdZ7mGsdYPPWN38/
ItRBnV0m5bBQcr+tIVP2wGI4/LLL2WrZhNFyWyaL/jqJhpUikebFgfky1IRlZWRc
kox4+26zJq4Upai3bO29KzNDdP+tU8NkmwGtTPtHE8NVI88/oNUW2zcuT6I4sWtL
EkmS3ehUW0NqSJ55NNbUqdjzC5YTHBv9xZycLr8qTaA06/CK//NHoau94tj1NmsN
JfLIUJR6mvPTwRwrEYWnOohZ2TebggK2SJpTYRasjSs46LYIpjcDn+V8dLsmfLwc
UpSGKMMMYtUVY11TG7UJVUYz7D1dRLs9/RaiCsdlbCT99OQf6tnU7IXxTpcqC+Y2
ELdI/9UEwqkR3ccejDIq9leob3D6xsL0wnQmQTn+in1EGb2ZTYPEuSazVk6P67mD
H8Oz+jyCbMJUo0j91xjVSWIl3s4mkH/SsN/lgCwM7x88QFJ4pexou6rFPcZFCHal
IcAqRVya1K09leEjw874cO5w5S5WgWgB7MDK2zfXjARYWPBrcaX45xkvDuspSt5k
8iPcMw5F3r6MRd2y2YJ16cX4tjgEL58eAh8WgtGx3BSYAJGzv3fXKR5G//ra3TM8
Dp2qNXL0P/I9nktiYarJaozQ/Ql1hUM2qEJelqBemmiSYlqAaH4WyCSCLi/NA/vJ
kg/UdD++Di2nQDIw/nR3KgTaJGJ+vqb7NvjbyxRQcr7Gxl4x1iJ4iqwo9/1rdrAP
Plr7XZa4k4cNT1Va3PVHlsOxq5dm7KHQ457nBehnUesNqS8LQyoKmKk3OqNsRkTA
EP6NUJBUSPBF0wAB3awMf1ZBk+zUB2Yr6UFdmjWIPFx+/1uhS+BxsETId6+Ry3Gk
Hm2YoGngqlrDrlQ+46Ta4/2OYHZuKkkrrwkwWjkg8yqVej94sT+cTxhB2eegIv0G
fE79+rh5KVHoS2oISLLiahIyqgHVnljab6LQbSsW3MHNUMVOs0Z5d8K4h8DPssgI
ChF2f1a++s59Da2Ty0uNNmH9N0i9d+R7IgRwpECvE2VW+d+ku2WQ1dwb2uiKsbL3
vQi+KjZziMB6R8FPSPsI9guruSwVHLm1QjIaPviQ8u1vNgokeWk4oLh6Sqs19szb
heclMFdUUJGltIFUrC5FV1Ek5hGJI6NhqzOBBhwulrYTJnAFfuOBMZXeG52OY8+4
eFZ5CVITf+SrXQbt52laUWCC5dDlTt+dW00CPNaFNiKR1qKV19N/Rc8y54YuIgP+
hPkASRhuakGObbn/CmAOBWA4ZedTWnkvEQBHJgZQc3Tjzu2BB5MO/nETlmauF4jX
keueV+jhDwuASOeJhhUTB/aclI2D5e+VPT/TsEEKx6SAdJA5FMVBAcxH7xuq20Pb
UbncwUhAfGGkr+J8nKTJx9dBiWbgNGA71ExX3yJeITXQPSAF8dtRQCSOOWswgffh
V3YdNjHEnDGsYbKhYSXR3NkbBzrzMKlZ/0DLTkm4Ga1TBpHOWWtLvn4MazSYpD/v
pHtGPY5SvdZ4mvrmCd++rHsKZmq8AnmT+OX4pzs1ypDjgrgJABJepOYMJEfa7FoJ
8USyBFNZnPf5cF+6Za6BvwK0HSGOH9KUmuX90jwso7yqp2vCS2unzN3//PtRKenb
CYbiIaWfvpU7d2Xu6l4NRKv4TZ85SJiFImku3J+HmaCTdT8QfQeDXTVySk94mvo3
iXsCjHiaLaxBvUvr1gpf+ovvJ3df6EzAylhaNFZ5ndxZCXs7/G2ysLlShgrCwjol
ThEKysjJPqGSoTKg9ESl001is3kchL3FM5CQYeosskeKed4oLb6RfqdjxtcuDXJ+
HIQ2/Ml3fl8eHY2m46O9R44B7/HhoCfpQkNdD0Lzr0/PMdIMbMML36IiWZfi1lmi
7YS37qUxAPYmCQdhT1BlVRi688BhJeVffclL9fO8dCvB1eC1TS2HTmZXVtXuX3ez
3rnnYSoHkp43OyfPDljHx4VeWmEuU/eoxlCmiJ72iIu8TeBfhTvZBZSMUYFfVi0Q
cUgr5HvGYmLZMXnV7D+qup+ejTCrTnP9eGrkkdnqY/PCHHsaOVxFo/68yAyXtfWA
OKhbkv9gWqn0CGzoMupZ5ILiUxKI5GZw4/X950oiXAldmOgujG+Dy662CzYvdMsX
uTUt7zZhxdUrgMhCBdRIb+mOb1msae+gtym1eJjxsqPWY45REePlFbruHQnX78W6
ybUHossyWtcBYevU40S3BdN4osMNDBJz6dBljv/JZNHrfGMzKeofuXawsUNTtdnq
bilF63Z+7NHUcwAwrHLn3u542s8Zj/QqqUF4DKhGmQpDmm1jVYJgsPr2I3fE4eGX
LH3H07npO7qhxsP9tB9qNF6X1ENVQjyUChtd7zYHKErR8Q1FNP5zEKbfeMFXsz53
sw3LYqci6Hl6CEjtSprb0HY83eS+qayGiGkODhaY06c1GJNylWiFaWKMYo+/dUJg
Z6pXzhTZWtEJy+UwImzS+7JE9a9lCm7CMmoWj2PkjKLFme5OfOiTKCvTqgs7Gqm/
ITVLeyup8anfs3R6nus7I2mNq4CPj8+MSHydiRNdOgIebmGCeS6MFivrI/5eh+jg
VLT6aj2/66K5AB4lg0YFsZZJXB8gtV9nzOTmN9UqCecFLLbiF0FfmU3uhURhQyKe
mlMMBZp94pHJu0oI9/my25lGIchyCvmzG6PhahnAQZ/es8fRvhID0gUeCQnNACSm
i51yQnuP3On1JXWdjpQ8e6f2qOtMEfqEUiMZy2xCTmWridYR0kYJovndeI5qvwBv
7ouDTcc/wNfWXll0HXt5uqo8pluhVELkRbrHBGgSGTZ6uYpbPPkgTblgJHoKycEJ
+9fTWDZWX+r1nPJZmu6dXh8+UShZQvnKyplqunO4AXlHqEF8jBEyYZSujWbfYJlh
izJaRqR9i5Wfz8A4PrudPp9GftbuncmE5W8os/pUn7GwqoU5Zswaw1NQ0wsr2snV
MiteHUwch/QwckDXyNNiwQmBL6JN8X1SD89cqTTWmyB3BzP5pRbQ/trc9Lk2cgmS
u1fV8P1C68fzZANwvFVl2CnkD2ENaM77JFY18KOuT1FznyOQKhLyWeE+q2wg/MwP
9hJz22ygdkH1LBubBib+5uV1DrPq2iy3iMDU7cI0loLklKIedXN0KV+xu5XyuVE6

//pragma protect end_data_block
//pragma protect digest_block
hxhLuvSHqj7wnD0nTarmWyON7uc=
//pragma protect end_digest_block
//pragma protect end_protected
