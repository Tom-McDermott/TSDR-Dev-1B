// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
sxGk1jipjLN61T1ff6MgvHmzXhlQtloddBOgerH/JgaIjdWnQNrhW0LL5JTwurFYv4WPH9ERNw6V
QKQyRl0mL8Zsg4zKXoLhOrYCWr34GeIiIb8s6cMrvV0fhczsugIoZRT3HURshDlxz3BkNev1Z6qD
+OaJqq5KjTEIXNCE7RMO8/tHtuWNyJejdVPspzdfrRjp8JLDRDiFNDtBEx+AIvdJ1FYAed3i3KHZ
5EhwbgIHhvd8cBqjQ80+PuXmty9ioZYaMTdWcjd8svu5t92PaumIFiuil04crnn16Cp49wyVFF0d
i5g/cfv+XXp+46DJg5pnHgY27Wm8on/1SRZPog==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6368)
fmPp2HTAZb8YZu8imzV8FlRTvxj6UOJyBhLha64hXlIw4xrTynb21B+4S2H9PJLs91v7uwQF0uX8
M2P7J/HZ57EhaqQJAbNFUcLPscW0DzTYu3hbgOpNKgQkO/8Q7ukgxquPGYT29C3zVBvuOL+lp0sK
JbFLiPz1Za7W+gc7q2Gl5U3H66NL5EJl0eDiU03tkEbatkMn8KJmHibINme/9oBYOUGEf07uLttQ
sq53NBbvGO7nJl0856FOY0JaRsSmMMKNfek/zunsI6nvEpZ+I/4+7nF2Af8HLitdONCXyYncl1UH
VnyC8JOvVw4ps5lSjA0tr9U10uBYtAr8eMv2JnIpWbjA7+nZLCe/taDyw76jtycoizFrwYd7dXDe
LZZrw/kvdWMivzaWm8gNWY1ul1vMhzMMfrlWx5mSVEAlE21iteiqy/zNmVTTx9yvjeJ5o5XxKRsP
sM61wpA7q5XV3dWoJouJksMkJ4h3SU6i1AzXgA2dwnv2yy9Q8DeZtnfbk3iUalpnPzjCKznVYe0N
XvZVrdGr/3Q/o3KdTKCpAkXnySJsYfa46+dXkOsLlsIH+EbHaWzh0wPsJ5oD/It6gRyNaDcEbKHm
ZXS9Wmz7cdUX4J6qjebP3QJyzTNNPK+cTpiigJgSAwTprBmuGAwvcrKkIJeKnHM3J8ORhCuZybK0
PQpaePAZjC2gZ2IyIW65wdCzP1mwkNXUpV4t6SR388xJMEZyQHFDGXerMVctlrtb1y40IHY5lc5M
4MfvZNlbDiSxC+Df6m7TAW0f+net93ydXnfXRd2YJ/UbMytfOQqlYgoXmwd7aIckaE0fCnYJl/gl
4kFArz0K2ClFeMsXm3uQQhR5U+jJ1udpyCc69x6wVjtHaJobZNM3ZGTn7UDmOUV2jxknf/NLvaU/
uP7kZsxgL0gb4d8P2KylZwqOsITW3wRc/1KoSrHjq+ymvAeNJaBu+eba3GK4bHWv4We3uEVNBcW5
yYlZrRL6nPZbUFRhIwo5fAqi1OizThdrBTcfiUB973zafAZZiUwWHoPnb1P3WypkIZjo9gQYBkz8
xn8ZjO4eMfV8KKvHMYlEUGJBb31Ss1PaGKCo/kXdprzfqNaRgm7lk3AbfArXuaDFlcQEF+bZ/TUD
R+URvbBNK8eqFyak5jC3GKzYcvBXiqn5utbpGm4B5cs9QY3WHHUAeTXu/LnkhejRa83QdrXzBFzA
PjZpqhVr0quh80McFmhvoWakmrN6HKD1K1mPz2iPpAD5m80LP/EMF0ihw9df+bKS5Oh1pa4MMaMK
f1RZodUF4Z1G6vhGRV7HiOei/C786eMXkPhU9B4WtPQ5Gek1VmeVZiWV2vYqK+tpE93GSJ/QmDsf
dDRwTJ1mBetQxblRmvaHAuI78PZ9jxNR/23HUcQKP7Pgba7SBDe/KMOAk9LXGJaL/TIRO+cds07a
1N9A6V/LsVxyFaOlbcBWnviLM0cq1XbA6Shac4HVskoqC4ynxxsnKmr5HETyJhfgeh0kL+I0l5KO
SIInYrR+8OIphmFLxTjueNDRKpgkwKfr0EEWH4gHZNTOX1rMAkZXu6LGC3fZ45uyTx00BbE2Vtw5
r5A3O0e21p/DxzMzOZZbA/b3etZwDhh74Vn+iey2b3JPQOd3kzp8zLv92Nf1zEmSvTeMpHplANmi
JAXvjVk+1YaQ5zhwhLNtB62jlmoOemvYGXmtcQy7o8bXjs1BX8zS2aWB7juX/sAKZMw7WqOXRNZE
QceD/aaFqb0STJEKRSUri6r1jhUQeq0Moj6gBSoukJOAayEy47qvS/WOucJeRGzL/ZqfA2+Qs9uD
5WIMU65UaA/t/tN//aH5ZQJWOlFY9+KNo6xqpl75K+xK+VVUExy+uPBxJXpgLGE37rasaUaq3tNq
M3mCv7wuQbywV+SxM663zMdd6HseYI5U10Lm94G5uoP263FtjjQdqoeDmfSY7/pJnvh1aAFigD4i
+n4bsNx1ZmQK/9QoNPCEz/LhUmf52a0iupleKmA0ukzHCOrOuBFe6Iz6owPXRwY08VS0murrQnah
WR0zOeFe3IPb/6WdcQq5k4mKdJ/H0OwEAd23jBLfhYpvoqtpZy613047skbcsdGvkLMh++/AHq53
fLhpYRBTHd6J4BvnBBB8m6UrAOHdFOFa5mh8KXsN+0tbjhOPgCouEMu1KlHcGeqmi1OLGVV1ELls
N6++5poIXw2+7jvXE4SeoWOcyKaapNbjHBnKde/S8xcgnozjl+i66j4qKsdh4FLXtdx8FkRkEVvu
MP4sa0QyKL3YcF2xC4AyGJkUn3fQ/BK1A6i7QVydAiMQbFMNH62lFQNmJR2ki7Xsww7S3uLo4IQI
YPVtv0ublFSWB4DwkOkSGilWQIRp1PAtp8nOgFyQuytoEoEhscKkz4gFjm9fjwcnBtp3oEDSEE25
jmjE1HZ91/gnWA1uH8L5rcEPnklvj8Kd7DIRd4ie225xwV2iJxPck8NIOVx9cdPTECsRJ/2NMfpB
bsEWr7N0ikfGDobBkHYr9ydvJr3LlhYLZpRaTD91+8qPeDNIedW0eVCRNdpJ1tKIeWsw2rBgr8JM
2Uty9wcWOGY08sGIjYhTQPu3QnhYybF+enptynDqJxQcXLRTxOOSGXx1KP3c0Rl5bdbvbZcf8pbT
l5B8A9/YsCPzveDO+1m24GbFq8UCq75r/GoidfwQYpxHDsFzReh4FTiQyYUlBaaT915B4wxNH16n
DrlrMaZgzPpAeeRMf9uSsqNAW7BLAOVZbJfoE98AffrVbH3RI7gdJell2BHqfXMsfBHAkIqI22sy
u4IusydoFwR/aoMb4qkeDqd1LNybutCaNnibpdN1/A2jp8jW2TSLdgYwHdLucxJvU18vClW+dVVF
RlwaJEwPiD6jgvWlMr6MALEhry58nXfdlpHUHiKIQe0BLMOqVb9zMbOdS3DIElA0lA/BcrcaYAVi
lS7hS4f90UzgFGekk2ZA8SQEqg9qf1U0K4woGtJUn02nffVQ0PimL2i9TWY4lsOqvwTnsdo9qshB
yjKiQKfMiu6grReQY8wZwfFVm30SpuXLSpctlqz5sTf5nChk6KlGpXrVuymDrN9YkNGvVK2CS1JY
kEmspJF0vTY3Q7fjEr14dj72M1rokxGqU/NSVSfJBKaq1W6LEDSXERB8Zk+zp1J2lR4Q7Buwd7JW
TZf3qk54LF6hmyTOuDVJ41XmyHzD7pKmMclvwLpJjCrl6wQ5Wlq3Y9eOCzKdxJNajtg5w6LEm8da
/kgx4MBtOHoh0Y90wAsoIDXb6TJX0vVjaJ0DtC2bT7F1qPyJiG0GuSknkfou+zvE7OfqcbNojY0q
gz8I861M4jKXCiFe7oyGJbHwP//nfd70uuKL+DY89/pbx+6OsVOfPgUcV6eJPKxby0O/sxfgfXYA
t+Lb3P9TjTihUhDFF3UhK1+YxxnTZMpaYWmtDJeqnG0s1F7XVbIyh8AODd32sEWt9QnCcXlsDiO0
930UdvjErg5Yulg41RF2YpNpCY7Rb/nzfzCIAiqPk5Gy2dIi6cM1ExuU0E9S6z14qg6kCro6+1kR
wjkyYm2xefBnFXi+16OtoHHD2MvHxAZ3uMtslJhTRsY1QbnlgE5yxx0yoBKKYUb6u7tShBvpxSxZ
QuRUoDYgmCI9/s1xZ1Iu8AwkKYz81VTraP3aea5IYzJoMW505SVMFfeEW54xY/vH/7fB3G7DaoZ1
JmHn1S9/xJFw66KqTx4K0JXqYAtD9G8irDrIvj/H0WecEt0thMCPt1a5IrW0+IMXcCq8yG4waT+4
5CmUuox17nTZ0vxaf8cNRTE40EgkhfILvEinP2p8GitbgDNJHHfq1BlphN91KfrlhziyiJvvUrkQ
VNlXKV7cbenW2q82WRW1wblQm43YmPhqmnrxdOdj1d5YWiJgFVMS6Z+/5pVu3w+4WjrxzRV5pVmX
XB9x9wqfwSlgWvo9epBqehv0v4dfyqyUij5ZwhhdiRundd0XIIo8tXtYegbNtK6LgulBxSYogYI6
qZs+ewxYBD1fhUrLFZZAHHCeRD5tfCBE49DHnrhio9lKN6ZopFhcK5P+sKJ68RV0cPcNwVVg0nK+
PIXmWXXnGimXAamPfX9MvKgZq1wFHypFhi5VaDZcf/nwi2BuqJeAqd2wZp3YESVuYNc6XAgxutK4
jcJCSDY25aT4X2EzdwURJqGlqzdlDbC58zJ+igydnR8osStBzTt82MiQG7mAT/dnGcSnsTsuTeOe
7PI43azVYpAn8WVcZLkIioywjfgWXPwHIjr6cq5UdS6bLtMnH93OhDTeEyu/ZwTxP9Vp/Jw/H+p+
zplLcvMAOXCka7YU4SV7U+xoLFSDdfFK+rBeuA5Qco8R7SG2iZq1J1Ah5f/jqUEsSQ0S2/BURuXH
HvkcHotyyWudzuDdqjspG7Ki/sU22gfh7iiujLAKKUVXvFgmhQV0Pq/l2a+fBkfpSm9DQcJ62Khz
oZ+Ws7j6T3/Cae992r0VyaHV5/257BIP8877vYrN6tnvmH1LaglhjdPJGxZGqASHaGIfiSd+4Qm3
48nCozD+PJ/LrbXzvx8We9c+0hXWVgYj11NjFe+bMhz4HSc5C+41o420wwOYswVrng3Iyc01UhXr
69F07FzGudX06GMl5klpd+Fszx3Q7MJ1EThC0EAFW1zOf/cH3Ft33LqNE4Wv2OOxQd/yGL/4p3iX
EPqfqMMRyVQ6EniAsdGVVvWLIzuUHHomxzqLzvV2eB4Q7DVcmgpAe+q66AHBsKqB2QV1snILr+cH
l3BPKszYboeszuPUF7qPDClvkTbXhxoq3OvS5K9z+s15T1TXYE3XnnRYhLZIxSFgwntnRCYzjLlw
u4ZasvlP16Spk7bsRJbXJskO/eGxp2NQMu7ZA7SELD2yW1AwE737yrh8cmJoTnQx3KXEnUbZ39Hi
bD3up+aJgBxtshlVgk6xpZw6cWdvouipZjTSvQY5XVpSrrTuQIG7+hm4rk/ewHaihMHK/xekhbH9
9GOwwb/bfo1iElOh6vSUrkJGqyeLomcFWgK1Uk+HXSyRs5BmoO256MGWtpxYkl0l8K4YY9gaHPp1
oYHW83gEsKc+YrF85yNnzQpd9GkgbGmw+yqvQ0RaAXBfUgW05wDaI/2aFX9/0kDrfWtHHFHjqN8H
bifBWaL39LUCAPjUtnBEZE5h9g1jX5iEvSaNh2MJl90GlQBNzWVxilDqnpvnURVH7+OqPhODVQ1Q
Andw3MwQkCGf/8ZYv3jdLkYccYsO1MBKCpDujXb66PD5K6jgsHcCBfvJxsrjrlNTJCtjLo6JMpea
TpDwsY7mUNkVyKSOK3e8xxu5AEZO6izRMkqMib36Zrj28O2J10cKkal/delE61JMrb1ifWTYitTT
2ikN9ThYPVJ9/XFargl+DvMkNS98cJh2ynismdMGllV+yvf23edLNsMhN2x63dHSTy+sHHRWw1Vt
CJhs2a4/I83iEIbFivAqLr0j3LmiaGKlHXsaOoqWqvZuTQZDRD9v5KgPS8CU8O6GvRf2xYXxhUxo
AqdqNyrUmusD51AdFVsUG10IPepdpF3xE+kVfv2bK5jUPem7Idq5K8CMdojAEJDhOKL1qOXdabsW
M5Iw+dlv9IpHGAiY/V3TTPK4Jvep4Ezl+9BoKKfsDfu5SPPR2xmMjTazUjG5har5wH40Jusme7pE
6Of+iQJEid1lEn7+dU/JYgkp/5G2v3p+FRfhYx2K87U1wkcTxSIulo3jVM3aSfFDkWFnFaesvt14
3Xqk5I+Z3qi2H4C01e+n4fZfXkraZhecKVxpsRRp/OMEf9HT+vtedQ9LUu+Qt378aPMvRnns/yf4
FaBk9mJhwbh2DFuhjTApGtTRZssrPkVyhQQbPyh6oHWExYAio/cKJWcfnfLCKucxzCziiPT50H3I
amiqFSxqvd8HohRO+4bevUrnOPJiYB9vzYEW6eigcRnfZyh5P6eh0JWKsI8FsQ2hhTcjKEMIlnBx
gxCRCBjAVPDf/BQ8mEgdwnaMWL7lbbiVc2yD9hDv8aIxgXlKnwJdPjVj4DjMToEet6aR/xXpfPCC
Dv94yGL402/oqoLmqtuOOGnKTJxPAFct6WxTPovx6N7oX/EkF8MZN1Yb7vgJCd5gJltQ+8yycP/B
yQiuoAFg2EdpntHS3bCDB5cMRAOk1/RlMQBigKjZ5EnQ4cCuIMdcj81oVUJcWUTz2peFWadFW/eQ
kNtZKTRY11B9Bz4nPxAv/uS2sxcxEj4BfWi1SSEtEBuB1j2F5o1LCSEZgqFJbHFMsvN9i7oTCBTf
ud6xXk2LGOtLY5tsWRN87bj7zMYwHH83iYY8S1gIP6O52/tMRftTGhW0kWyna/OPbh7kSNcUc1NX
cdQUgKJ+ck3aRgN9l9fWyx7Ru+Oh8DwH53VOeWp64pNn8J8vl5UL2UaBE2UUIqgwhPlu/Idrx/T9
iP4TjWq2zswFEuqh+vyFXau524eLauAFjdxWWTF4StkuUelhrUbVTQof15mxrhZUZ97vxuYYYvnw
aCObe7Ti08R46pF5hZ7thM+lF8NZLY2RolATLaAFlZ44WnwJrzItNFWN5Hl2gRTrZkTQofVXdJlM
t5MK8BvY82Uj3vEGVmh1uk+N9HGA3l/izm9LZvP9GT93AfKlYATsK7c5CW+XjGZDqBTL4ioSTvYs
qSptVgl2eR64WS8CymKeYxXJDDU7LYgfk5ornAIEp/oaPWJ7xnIn5mgJdpuWN6nVqpXS+gjTwsij
XHXab/bzU7B5aAoWa40FFo7Zoqcq+9ENMAZV2Js/A69M48LAtPA0Y+BtzDtSueMw3EqLyeHlo64F
IisjUTeiazP5oqMwrkoFR4CPmcUErYYWkBLrWGgsZbji/auhYQmW9N/GQmVTPN3gAsOLw7w0m+3l
lQVIcY/YgFU5rqX1PmZQ9PREh5b/OSe0UwgN0b/kLnzWhA4TbalLZ3PhHMaym3dGPZim44SmX1QT
0+btawS/75EFtWM64b0iXnLZ31xPs85tmhVttcst1sHgEgnWIUJ7OS88fNUQANw11TgrPCeQ+vp5
g+WK5OVr2OGk6pxP+qLfaHqH/1y36angXdgFUbSsp6eZlMJqKHrga/1A9Ou0rO626xgNvJtT8rhc
RutfRAyDs2renSQNeotmehwHjVoCQr3IoLF1Iutugjiix6EkzouU66tXevR6Ty7ykguJgc/56Pqz
rUA5iqJVXLQvOTOUrwgS/8mpg8+lQCtCSGOIXm28OGLYeiovFKyTOIkR6N1soUmkGfZ2+ww0peFQ
OanM134/3iGuuwMLcqhmNdb2SmC5uRvWSAX7nEPM/gXswJ1lYlHUjbJwrgXISjQfzqgRNcY99zqh
+XlLEx+q6VyVk6dhtEoWNqvOztxt+OxLxi86jZn0H1zfmN4M7eU2EY7SPvUUTTkWsyYF1BlePOZU
+ecwsK0XQ71jra1qlIqWOhjVkpIeVTMbEPilg2skRJqI266FU8WEZnHfuAv7ZikoPv7oGnZFSi7P
fxpbRb3KxR4Ld7FeO+8bkWbvMV5qbAHJ+ddTCvgdYn4mOE9+ow7HsoPn81h8dmG8dIqMJ4ZKAf4r
t43AyE8Dn1L5OXR72jNZe7/d6n4+dTiK57Z/wzkTMYhr+JiEvb/HgB+yzTGs+hrzm3P6RawaH5LM
A8BRmqrZZvudifNIlsL8MwvxlncRZFOfTb6zwt2/FQ+dkAICyoRPi8DcL8QOit0HGcdU8D7y7BK6
W5a+oZJ81W3FtBDYg7bMdAlyjZ09epTphMGdOb5CjuHW/fXXglE5hUl80GslNrMNaJKWHYimFWLL
+wjjZl3/k8ZSv1/oaA24FLEvbrRTsETKTZ5U+1qsWIpyZs1/K4OGD2ESbB+2n2PcVmr5HalhQE7X
PgWZI7bg+hpKgUsbshefJOkcyckdF5BQPGRTBi2obWy5Uh89kiIxXXuw0Z4yRNL0E0TZBfKRbf2f
N8ZjjfDIYfQ7YCHbdRRwn8yZF651DICp5jI5Flp0dPrRKfJpEibLnmBi5wXvWINneub7iQ9WqTXi
yZqETuAgIj6GUmHLNlj4IrGweRhpJU4+wTXC/ugIjYfF03xyaxI9zr4GA5ECdx/HEA2d8bQBwu4I
hQLDkZnYc5xwRYVCNI80Tmu2+fzxc6PpmuEgvVTjx0GALRuho2xJIgju8gHuNB2fs93Iomvk6paV
htBomdCfnuE3HAVuU0rrUGtBD5AkhSO1vn4hTGCYHxDpCsrVdAbEY0oYoOTGvqP1juQshxkMorrt
JTeohlFD/U/tRslTQcthMl+ylkiYGVSMoyTArRoQAkFcVeguD8uzpAXenUBp4/HVlinZ7ekYQuic
L1ZhoO4tZYdNVehSKTWvWJ88yx+p4hxJSaZIPVAZy7817bktMroDu/GEJVVdK5YInCN3CYJZTzGu
r4Dbrcn2UmSbN4PvIFVUJP40Qs/ghLmIrsC3hLISicC61x4VO6WHgUY=
`pragma protect end_protected
