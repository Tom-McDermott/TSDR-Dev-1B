��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D�����WUP͟B~�ㄗ�g�:���e���%�)�R-�{%Ƕ#�Wc�Zld�n+?X&w4
���c�t;V���?�,'M:�rC��cB�o9� /n6f��0�*�#c ��p6��JzR( p���Y���&f]�Nƕ����oΊP�z۶����\���r�Eg���tt=i�.�"��i3Q�8��^�|H�0�?��ݩY�4Ժ���9�W�#�H��Ĵ�����qSE���y1/����z�"��> J�"5<���ȟ����,<^��mrq#`ހ~Fz\n�T7C;��@g!����ޑI0(j\Xx���U,s��z�������Bs��H��A�w
�A[�4�zZJU��������F{����~$�p�FJQx�:����Y����z�q�4.t_���>���ވ����(u�V�"�A�7�FA:����s�^��D\�+	ݤq����r���������21c\�\��
.j�� h�vX�D�X-9�����|'nmp���B�����#N�ķI����H��G-b]c��A��H�0*ο���w�]����r1�����>�p#L���/�A�j�fU��Y�i}z�vv������FВ�Q���C��6�bZj���b�O>��Z���"�O��Y�32����vMq��ݹr��:��[����.��\�M����pk��}$6��&��e�>~��_�^�	������$V!X�4{�x�8�=Ds,�v0�P��8�T�P�]Ơ�m��P��R�%�A�Tf�/�Q	�p�Y�v��P�P���52xS��Mt�>T�W������om�zP�l�()V[AG��D:*+���w���<�~��za��y����h����9lk�^D:z���B1��Zj3����|]�X�H��`ؖ��V��t��-[��S�<h4N]�|39���m�Q�x��#�o��p�I7�
��'���o%���̳�;v��*� 7�e�� K���b��2���Y���JO��< V�Í��C��F� I�z��%�[�/[�g��Uo@�2����#�})��� �a#F�w���=�]G��[_q�[��'co4+�B�~;�l���.7a3��7�Vb1,E ���l�
{�c���p���Sr泛Ur�*tQ*����hk�|�� �~u*��<�`��	�]�P�jO�Dh;.��������za�u>ȇ��k����s)!(�é���������Ї;�B�������P0�t��:��`":�	�m�i ��0߬,���
����Sy)Y*��y^�ؔ�'�I��&V��Zs[�d;�K*[wi+����e!����	t�Ł
6�rZc�sE5�TK0T�\��Vr�V%1�1a���;�k�KaE������L���[��J�h:�ј��������Q?���e?��5?v�$�$���:�EIZ��x��Q>�B�=�o}�]��>㑶��W��J�?a�&�*�I����r{n���e�dݖ�&�}z��`���r�+4W	�ۛ���{,.��R��H�A��'e�Qy��c���>���e���.��#��l Ugvg6�1TB	n	'^%��7~����,���q^�P�����
Hh/�ΔΪJ�C����kx pV�ג ��}�8/�B��Q����SKQ���J&��Y�h_J�Z��͢�F#�n���8���[p�z�ݕ۟�gV�7��;�DQ��g�� �{������U�+���ߐ��f�o��mc�s�J}�e��K_~GfGj��g��sn���IC#����ECq]r�:B*�&�>�˦`I>��MO���y��hM=i�M����R�f��n�2��E���#�j'�ė&J�+W�˵��^��--'t��a�k �P�4��_N�鎚)���$����l�1��(TU-�\1.����o���,.�����MS*�gO����`옰�4
͢���x�j���X\�9�M��lZ
��p#"-����]-�eV�0N��=Z��w`�@�|������5~�@V�g^l���b�!�&����)�y��zq�0n�9�*i���^��'�O�]�id��K� #��}���q���6�d�Oj��峴ּ軍8����6G˿GW@� e4se�s����֏���3��"���i���; x�M�\�N���^����AI��Ra~ih_Iu޲�y�o�V��/[��~/�U�9O'}شpIp�6�S6�jЋ��Ld���S�wka_�%�\����O�Gwyv��n3)�C1�QA �NX��^i����od$�S�mi����iDx��~�YB6��tv N��e+A�C66!��^�#Q|=2�^}�v�#]>�q�rǣ�i=cA$��,wW@���U�f���._�7�/q�J�"w��p2��[ߔ�:M��\�ro:�o��ePUSPA5;ʳ�\-��),Zn��a�!�6�<�JK�:C�R��M��\�c��{8�q�B����L�D�}�9��x��S\�8�&��@/í��/4T"_f�^�)�TE��☔��n~	7��6�;�$���I]���u*(A�%(��� ?R]��DXgD�#@���o�Kjي�۶��@�4	�c\��@EI=�뀗���f�A1�b�/ׁ�)�ؠ� �l���s����&(Z�et�n��� Ձ��K)}a�;1)�<$q�M���,4��Oʐ�w�ь��a�=�`�\ I����K�/�C;G��(��k�=��6��'գ5�KF�v���Lg�PaH���p�-�11������>o�.a�����;�?��Rg�b����ݷcT�U���r����\�)����on�'�/�dcк��ہ$:P�$�a�J��q.
u�B	�ۙ����5�4��z�L�ם����?2u4K��.������}���8�-�U�Ë��31Xi�`M]z��)�����B� ��b���gA2��<:`Bg"�bY�x���D������>��u���{Лω�
XB�T�Y͌��:VƇ����#6[׻���<�'Hw7�,��X��g��u_����XojG�S#mT8K��$
�'6e�O�]�R�uF��?p���k��.m��;�1�z&]�/����[����?��ܥA5���QTY蠰�yY����Ѭ�1��Э��'��3�d?��
Z�»�[�����}�N1��dQA"m]mu�����&Y�(F̈́Զߚ�,܆RZ���-�ښQ����ɡi�@~���k��x���Ϭ�(02���t]y�0`��4�+}I�y3����O���6����i��ۤt�a�[@�lN�S�yT &JY���(�t�'�g'���*̆W���Q�4r��wf�N+B��^C�1=3�j%ۯ]]wJ �>�VW�f��&������,7�1.a_��\�F ���F����`�폼�@0�VC@��6����ד5ˀ6���Id���m����c�汅|̌%�N���R� }��yY+�2Ih�!�|������������Os� �VM�z�U�\m��زun5��+$�yW�Y0W���IG�8?Etd:a+O�6��˘3�@��֔/ޔD����3!q��~�n�@��=@����v�;7�M�FF�}֝;9EA�jr�B��2����e� �&V:��JPe�KL�ؙ��d�M_�1-E�'�f���z��v/⃎]�w���i[�@C���U����n�<��!{˃�+�J��Iݾ�{�?��B��H/��8(�3�&��z�刊T�6Z9�:b\x�R���p���M�tKe���VT�rcV�V�(�"��ye2���"G Z=j@�MEڸ1�+� ���W"rԉ_�[�A� ��Z僭c��n6WӜ�:PZ�gH??����rU`��O����2�/`2R� �>;�7Lprٱ��ET��<�r(0����3f�GO�[M*��q���,	J�t��^KB�FK�>��Q7�S�b8�h�MR����x�5B�\���kKsSO;��K�x{$�?11�o�-� ���cPEA�6����J7bi�qs1�0��T8��Hf���n����C�߄��Ó��d��sw������}Q��Ȗ�p�f��2/����PqZ��D�8��P���_�c�I����D�
�W�Y�|"����gJ@Ƅan�a�Z�Q<����~ z��a��ek� Tƺ��}FX�uqT磡�U�^{��A���=�t���vF��Ka���s먅�6
*�h_=�B� h�Q��� �uTd�������š,���[X���I���{�1���'�������ft�n�'��aRsa�t��?Hv�%�^��|B�p�ح��* S�'�����*P!sT$�����g=���u(IS�������$�䕪�7�*1�fv��
�l�@h�?������0�q�(/��v,�(@mPF�x'��g��=�-#�%��&k�Gi���S|�7lT篰�d���-6��//���
��x0p�����f�=�%�7��_�\�ls�/�����*W)�%�V0��(Nʠ�!�v�)�`U��u��!61V+P�R�3�oC���obt�4�,Y�y*��?��>Kҵ�N�΃�6���[��{�n�]K��<�V]+�0�����z��TW$ɾ	B"v�Dbf>��ozͥ�I�3��	��+y���D���}5(ly���2c��G��aRQPA�$��h����~�N�gT�_*�<��X֠�Aҽ�Kn�qh�߄u���0�4j�K�B��G'���h�M��A�C��Q#���d|v��7�@i���&�V�Yg�Ԣ��:��iK9Ў� ��� T��N�ّ�xu�#�z��2�P�7t��4)c�P�au��	��ld.�ſ�K`�+�~j��]��֔����['3"�ߖ�4�����t��9�ekw��X�O�S������\�U@���Y�r*����ph$��'��+�w��CU]��!��i��񥕮�A��k���z��<	���3�b��P�"�R�@��\�<Ո����y?Jo�r�U$��<{5ç0�:I��~n�7:�g�<s{�ɩ��'����G�T��~uW��Oaj�Wژ`� ���N�վ��R7�1�H�>�S�EP``q�4l��ut��Hz�$�LTG��My���pB�e�'���(u�!��� �u.z��bl̋�� ���˛��L)���m������7<�`1��l��S�I�4�Q�Uq]<�Ea�ZA˓;��k��pu�l�P'f�Hqf�Z1V���-ţ*�7Գf2�����?ap+�cq�_1S	B"*��-;4Y��"F�O>���h�A��gF me��Z!���ca�,��y�2���wnm�D-���pmU�sP�K���
�BI~
B^��@�fĴ7.�=�ހ\��>��LTՐ3'Z��-"��������8^�RjW�qs֕u� T�j���= Ť��sY����]