// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
KC1wKPRyGv/87BaEPPo2IVoyVPR6XGEh+qEVlmr59iV83FvHTLgCB/IhM3uE0EegtOBtU4Fm3CX0
ppE0Ilz9r080VCyuz1rfi1AUUalBC8o2XZEmnraFvqZuLxYfG5FHA8rnOFqktvvDFBjpYDaWwN3i
NwK5eMWD3HMmFrT/watIHSgczKXmLMLIknVUBnfD0w4IjvpPjW6pLdXPkG/J2RJmR+b+ilu5bOgo
/M4ir+N5KWiq+afIO7HtTiTDEnQ1ZXEmhgObfAFnFi6rRpTfRFCuSatKWVHzg/xqJnvlIoKlpnCw
UNl6Abia2meYHv4O/qdmzqxjg7tCo0u3htSwcA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5600)
fghJ77IeuoYNcEMpjxZNA8GefUOtB1Y/0r7lz5mYpsFJ5zjUdk8Il5OtdLKIzAVaWVAMFXLN0rh/
S0gC7A60dOjFQRtsLVTTQXdJrmNhyvSv8cM+vqkk96CeI4rW/UCNqiRsytAuhfIgXbUY5bbg+kmz
Lab9YSKjmuXIrMqij6Rs2Qpvph9ghy3zOUj2jNKlnc47JNeT/EjC5f1hGRPyPHdcTnyEPXSiKtoQ
x7cp/FmniPGTJg6pD5UVONOIMm3YKTKswE1foFzHvwMWUaFHewjQ61BmJv4I47YhqtoRsfpg0cjY
mKV1oKWLHGDAVYCl9a8ZxeYxmTSs6agZHiT8Qr+iHUN03CjXiztDKsT40bTJ48MMtw0/HIendmL1
/tX4z8v0xmdHAb8zunsrfiQQxaLfBtd7VIX+FQHdYBYqa/DltTknWs9TZZ36F5o9fmY33Cpz4hKW
w1z1WDhTIQEv2UO15HCSCxGN2nBru9PB2eb2KT8sO9ULbMFZeyOxAoRM2ZiNWbAOpQpHDFXlfPYJ
UM/sT/rO+bKmwP1JVgocnW7d4q/banSAYDT3fpWMebMQe/QrgHq3n32DMC5NgLWwhzKfSqUfpgcN
OBxfuSbGYl9i7scvRau+7BOinGaXZDCRv5fKVDim3KUYCZXxMp7bTe7Bx53/EJOgC+oD1vPZO0IM
degUdy2k2U2UPfm4yv/c8rtxoVbo8E3ATVrb97/Lpoe1KF8RzD8+4EYPT+BbPY3psDmQVmQt/ZP+
Hb4wtMKLRXJsbG9PpUEIOugHGJblp9WJ+XX7AeyG8K/jr/fjcLX7Z/vqPevykJvgt6MX/dqJPt1Q
mtAVoCYpXiRh4t2roHnFwStUxoTkpJWz6HJ9nK3TcAZ8HdocaR7EYfgyN7VzUqMg7338mQVeSuw9
p+vSJvJZQiyRsYZo0NqgjCml06S8Lzyt23EjMDkt+/VGHRUgrO/wD7fqT50SClgaO63SGthdievn
+i/ZCZ7Q5zj0M9G/lQYLQIG7RcUQVJNZrkdT009BHtMWVmuae0P68DZaB4xgAy+HTD7G+T1wByHC
Q0iSxy9f9rVwNyTyDEnpw9dYf5xLr9lQAVlP9lBlsq2sIR6QsrVyRDQVxL6D6mlivA4Cj8M518vG
njdlyy2WDgSeSG9SnjRSUT2tlOko+evH3svSkeh8TVyvxfhugelsc8TjA0gU4hfpWmAFD9TWG4db
+WGY7dU+bHJFx84JVCpjVnZCL3mhSuHbrGhWT3Ir1mLer0nQhp7kQI6PnsihsXgdXzOeKwx4YAvt
+Pss3l5KuDaZoq69ylnvJTVZsOKjkPIoST1V5nl3UA1G80Zi2w/yLUSIHZ/bPVuib6MQcIQdO+Pb
39Ewof5gmI9zgWBJU92QfFqKNX6BBakKdtBPOZcPiQwT8tqGLRkflq3cn80rQr1Y8J+xAGj1wsa3
r6qdtgy2Gk8ztIHEVhAcT2ie4jr5zBNp71t/PoFf1SU9iVLHlVDqWoiFoMjYFk7dlqkIeT8fJJFU
ogo2eUcxnhAgQ09PhwPuknA57bszRBK8RsWTZD4suPNozpBD8DyAWDfIo+UxYmCpKieg+9qOKECs
/OQn7Z4XtJC8jaUx7F2xKmnO78pLW/WM9/uxgGA7HQjhcl9ikdz07q7WBmfcB2yQ4MJ+QUey/I03
351xUNQlPeUzzastcm3oR8PFoCByJspWH2ljRYbvO6lWrsNP1wfqwbtjeo+cNiM7optkBZtjRkTn
JcwB767syq77z/gIkKzzPk2CYayNHL29S1gDb70bBBEIwhDg6Ay3stYBEJ58PVA9I81HQ1T96joA
/Zo5eNc2dC79x3xtn2gWxpBYSb4Pxcdm5nrttH/FEj3JPiumENyTz2OE84fgDQSOY3CSFvsIIlBT
s7ZrBNobV5yTf0uKGVHVS7x6GqYouPk6cvEZg6iieIWIIxSX03CWdnYa4Cc09F/BXuc2SI2aMfRS
z+rb05z1apXUr6qr4Y8jEYQxx/WjL+NARe0FeNBNEMSKKcFOId2ame7NeGpYnv3OQw8+o3CT+9SY
Lpg4yR9mGq17sOtqIE4vO3k3pYxpIp9j5/Kfo+ZiC3dL8QcDPC8rYO+Ztudh4U+yxbR2hPfdt5Br
OAu+Nv24BaaFydC7ij1qZWUyRLfHnqVVSGSpGzIsmaFkZtNpjjcsXrpIIVjjg6ObDVyYoyYq1XLS
I1Bt8RRAQoECgVWldKpSCBlfVSi3FihhV1qq8H/HCtYAG6GGQdGxHyucyZZHUijHiQ8E68L5cbIC
LlpRMl0hGVVUtiIc9Vl6xEkDMbIO+PYgSdoIfjXuIuDWUftDZh/dCSlN9N216IYogXmOj5QZkOb7
RIgZDTGAVhdGYcl8JuEfhL5kUjI2n2HBAPEkkOzdBYPcwqkGTdfshVfcFX1/1nywM/uif/roRYQ+
AfZvwVQAikTSrBAcASQtr2tl+jXAqS+OWeAV3QlgeE9PI+GCFcJinuiYPvygY7vwsoQBEaf5UnBL
YnBNBGj5YQmMLuFBNQ+jngz8VIVKIQKy/cpLW14DsIkfBMDtKfDAZgxcxUFG43zAlzh0sBVcEyZE
ERbTX3RRZTm7P6r0uR0XNwjpsJYah/G+C/9Mc8RaqAQKXjZ9TQaZ7eLMMRhsG+5wY6dBgg+xgY+L
w3JgEtxvb+pT2o6jZZu5acBLE+5vS/QSDSBf6vHulWFEXPMkkPtaXL0ErXOmxd/u5ssWX9L78G5k
pvxPsYbbtoj1cYCUmdsymHszxSSqMwc6nSt+fe6F7/CyaODehGwXA1SJ13OFQHlGJQ6sh3ymFreP
IGItdsVRPKw++ZYlcahHQ8isAy6VJszKFhkwojoqn68PIt+cW1YHTx3nah3WBQOKiBo8tP+usrC2
/Rg681jC83MOs5g+IgTnUZ6wEjq18daRv5WSm2gEVnEbWJwAhhGmPJCmAubbfaWXRljlWd9Cenjw
FlbfoQNhHBWU826nbE2+QO7/dOzOIGe80oHWMImO3nSTEKNrMMeEa84cFfkwOOcA6wFhm9LOuuVi
nlhVa26YOIU7TlsAZy8Xoby9S+fz3/EkJn2nTw0qQGWis/FKitgC80mpYddgqJsESUc5L0ILle5q
atsx0rvy2yFhHA4hMO888dwZU44Kz+ujAuJmvvprxNVPH9+LAq9+nUHjKnBHrNOG6bJAeqwnmgxQ
/yzV2CvrnvIjdjMw4Q9TYGRNCFMYXD6uGYFuRe2e1wQK3dGmelaT5vI13va8RVWLU5udZNYrJw0U
17A2ZXmLmqEKFVj/oxNrNhydGOOQz/ZKgGJ96g3WR9DeBQWaQyl4Efi75vBWChRIFm++IHnOyTNY
87ASvt165RiqwCOA9kjzPEYdmI+n2kQB/KYm2D/T2QkSE5c2JOapMRiTv2OWQ5dTqtLFC+b8MYgU
EH1pVeT6oGOw77kcT/G/rV4NCpK2/Z3rN4isSMTgeSsKsX/y2ae23O3JBmF9J5oHrxjQrde81iau
9lxTYYno37ZLeCd5qpghMkD+SysXTezV13tOo9zPkBRRn4PEAzsvbGk7zuWplMVBnBdzm7O/xjPA
KaUZH9j2PJdsSgjtZrrHfSWw0BgogWVWuAJh5qNfA92tlG1xTJaVUjZYeGAxxfhZJm3NXpZ27B3m
H9RvH/lnCpFshtvzFBuVaUQdyKxC3fVivqq9pNmKGY/eyqOXC9k6hJyAGAXtDnU4ogL3UjR3CmYx
a28NDsGKIxjgKVG1Oo8G2wjKT+31uPT+zibcpAeIiC3+csdDa9QknEA49y+/52ToWD2+j/fd916i
7XWS/Nn4QlFyUSkL961Ulr7icrER+HXF/kl+HYFA6YGGdIrIUxBkB0vDWHSmWlgZnt/BpE7J4TWx
Dabmv+6XqNsUOUl987vyU9PDAz61wDrIM5h0Thej9UGlTisZCaos3AlXqKa9TnSriHPcqE0gv1uE
Cyv8CvuFgf7SB0q9xubPIT+QXOuNbKqnXnsCivNAKlPEH/+7+d09viHGzUa4/Zep2BDNW+5KqZdi
kffeSeUO9qcOXnjGR2yMIk4m2XTrfnEHjB5/b9dBtAWJ59XwTVXUapkk675u9nHfIqdlQ1bODyX/
k+O4V3O9siUiiAnr+tS6bBL3Y6zEYbp+cQE90J5TXs/mwXSurZBkQI3YlyJL0HNskZlmifa7v08f
ei7ZwMtlmNgTHRBcjqLP2L+Tk6hYphblyR10rtoqE8LiB9EKpny5d1ga7kuLoO4PpLazWqxfNKxO
f81lMIcD6aOXq/1TAyR3IeAnjJYlpRSB4V1ECvCj7jZlN0KzDjwOmvRrmNy7Z96L4+SR8I/6UJCX
WGvGO/RRXDfVhUC74ZHynvGKl3HzZc7durdry9FRLUMKtHlJvsP6ogTJ9myusQFy1XEX6mbIg/Yy
khj1TYCHGhD3FgDP8yHLasTtF4HTCPKfWM07gcOtxwFN+3Do0ynhV2AkBOi/BG/D0547dzaoQ6Qr
s+VQyG2YGcwLVNAQ3yEdUqEliD4zuVDCpLXq6iccJDEq8PdsLc7a3vY37NR4bexpqF5qyoZ7P1zn
P2WUg+aUzDx0jpkzfR1hQfTvFfWdVKcxMZbkGGk5g1bCEobZbWb2BGhswN9GwTyDXFG4Y3DpF85h
QGkUEPHXWQShXJHBzDW3vJQ2LB/RPqMIp4AS32Oo84KkMigz5yFVctEC5hpI8wbcnqs7eiSTcegF
JnIPCYKoO9677S4yUpup7BwsHF2qzH13WnhpNS9ohsxpx1p/sAnEYu5f0Kkn5twP/Y70kG1hdY4B
4UpB0GczV+zPIhv5C2fS+mD2YTxNvs7bup4bJAX7kNRF3sOV/0oTyphK2S+8kQTd65J2wOzXihhf
Xb5UU6udkqPgb+Y4P1VMuN5sRYukMGAoSYphzh9D/e7a9UXgnfsOZmJgf2Ho9hzmmenLLXJ/lOta
CD9pc7DmWaQr3jugIxV6UxMxWgP8XuvgjBW6XbX7CVV4lqPUZ8EC0MaloIMlLPqwPlO2zEIo6GZf
HBOBpf08UUTkge/6Cbo0R/kJRowo024XVNEXAl80OYj7UNc7K9lZOQaIziOGAL4omrlK0rf1Aa43
m/bvuZZ7T3w4N+FSfAfjh5NY7q5OIH9f1vDDT2ENBRmdP/QANW4HdjS1gswKS/TEmbkPhpKF9xSa
++pTo4XHTRel+ihIPbFuWrNGHjFH2vo5Ha0KCvRd0Ld/qe6Tcb6HZaraOR6K53WDUhaF4OzTICtP
7IkYr6VCZmwfUoBszRmWgckYzA6kIrv3wM5zXXvt0EatrJ/5AESawRFyUEmU0OYVWcOXfE8XX/08
dpWS0QbIbdzePfIhu/ty/KRXEcVdIDfdGBwBsg/K/8ixE3lvXpvwpAH9NMbtgdjUt5u3b9ZfDcLn
lTJIsDC/2Q/F9D+GWAdyyalpCJUCsMrl4brJ6IfOwL+tchYpOQygYTKevPj0eFgIfaOL4T4F28hB
sBzIggUUIwlAnsMhyZG09CHM1m5ogu4Jid2EbIMaKlAv4DqDOTrdY68LoUlSHTg3C6q+vLXGQeQu
UCwsp3GrNec9u/7nsC0EDy4G+8c/LPrFDlXhDInH6ch1YOUasKf8M+S50Hnkqm1OYKmn2N60ImTY
y7qrmOJ6T8sFe+nqqJMcuRbiUlQvAEPhc1M6KON8ZbUOYDCz48nTlGbS9I1ra/Gwc1Eeju550AQ/
Ln+jsSy2monFKv7eb3xVwrLK+TgnEJY3rEN7pE9KClW+7LHkOpBLaXiw+VSTYBGple1zVOlUSRXN
wF+LilshXtm9YzPhX5o8fvJOwsHDJ1yl8YD0//kTJQwy0IxJoD7WW960v3GxQvU+b5p3G6gTg6yY
PYtZz11kOXuuuQS2FhwzvSw6fAoX65ikpehRz/GcMAskWl0g1kRvE9Bb+I8DlsKMTUanVPWcvf3q
Ij49G+3pu1/7gQ6QUbcGnBc27KB6Ilzzx5A/ukjGTztTC3qmaCN1DYP2fCN73/McPxt0t+Xa4WFe
kw1NJ8Ns5cnlJ50yVVcgU96u4OqdR0T2+28C27+VYS+rsuBtPAgTDKxEMCj74NuNQ8Uf5VNLAX9D
ghY5Hje+8nYJpH9cqD1LKkLx6xyaW8UW/ADQ/ukXzNBVQyi1iN4/Qbr6vARbq7YfL3PlU2dqLk1e
tjJbXfl/si6q6bdVaCFfkuRfTx8nkQ96C+bpn3W4qjo8io30IWhjzP95N6OxfuYoCPoBnlaxZ1x1
HW/23RdVD6q7dYMImfb3AujCxkIdSNiI/nntw2RU7mrG8EbP6iqbdN3DIClDydCNvnkZsUUkPjse
7DFPS56/XpDY7jbg3lf7w6wHnb/dkDsc0pv62jD1Wp75vAhUD69DfWyqQEF+ftGVhJbpRrQNPZk5
Arn2NC4p98sjMdUBzC8ZScowP9meFxptW2ft9KNBo07iP/3U8VJkKARn5uT4rI8d9GvSbNP6M9RL
nuZlV4yRZdEQ1C3ZeuCvguJGyKZzzqiHnfhbCfHHkbC9DzPwgNcNkj+8CnGbbs1b9jkOx0Ilwxxh
c8wIEPZ8LS95RmjjUly7z1G1HujtqbfFMi+3X+ETFDOqgOFnRmomeulQkKzhu+sl3wOwAmzsGDZS
UzA8qO3wcN/clPIkPHJ2C4ozjQJCtvZkC4Lk6vxtYd2M9Xc5cJm2PzjTeG6bsTgtaDkhFYlXs2Gu
HFb4/n09nhB6jvxbdTQR1lZoStgPxNUDZKl4xUycHXxY56CnHBccNRRM1lU26tEG1sA3FCWPI2+3
bjd5PcZ/s6cdJiMjrZtzDFVVzYsRfljKlsGaA9vTk1fsVNrtPFg2Pz0v5LndhWRaamY4yvAWlIjk
kaEzHV0Ek//CeCT6BV26+bbJtfeJIeZ/Lg4v5URGaIY40WiMxiR3Wxh2SzTIDm5GQhW2vNIWY3Qj
1XLS4XIN/NkbbBBDJdsuTzLs8xtEMK8coghTX3uS/4FVNsFD83SpyLwuhXS9is5gCFYsmoyYdLZs
7DrsBj8WlSlpFLfLlmeaD1YG1uG1Jyug3kx8TRXdbVUqf9GXaOA8JwEbhdWLet/5FeNwH7BUxKiw
st5JwCRwBLYIVSRaPC20s3H4Tq7pe3eWmRhYFB03moOnfLw8wp1ZWPkVo2OSnayMXF0HyaokgL3l
SEePdixnynk8WKFOfz7lm3TePm5s/sBbcx+0Qydl4cI31v8w3V9lEjdUQQJLAgpOp6pr9i51xaEP
1zWg0bLH6dIrMx+5HLcxYVMPBD7hFmyMcqJwVA7c3dVNuN1El/tXHaEfWRe/wyUjYTpB07gTz12n
xjKjKwkohRWDq4PsiZMtLdDMKaYaIsfpZq1GQ/hZQbwdx7hG5hsj/R6tR/CMbBkuIAFOUvyQJ4I3
n+I8YGRYDCyfwDyKYuz1UPsJ+oZ4r7uvW19leqtDuT/LiwEy4drvhPLvKsH8aFTadntM/+AnzM4u
F8knq9b52zQI5dYwOd0=
`pragma protect end_protected
