// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HFF+N+;CY):A1B=LK"UQR'L0TX8$Q20VUVH7I1_B#QG/0T?)D1FW#P@  
HI7#O)D1);5>>KO*1 60.4<:0HR2N"*@L#C-"1[+.'^4.('[WE GFIP  
HIK$SEY0[7*N=L6S#1IA\8NAXSVQKYZ- <8IW,HV=EX&[E%WZZA]@B   
H(=514H*MA]LD$QX%D/[%G60YN1PAE"%^@<0E5_ /KNMLK((;SBUDU@  
HI+&EP=H5D;PI#^$5G\Q/^@0=.0'@P;SI : ?F.OPDQ60_;J46I>2@@  
`pragma protect encoding=(enctype="uuencode",bytes=3728        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@U+&&S/&!):XQI'&;"F8XK]^;VS[&Z%[_<(Q!]\T+OS8 
@DEV5ID2"(H.=>5^,T6[4U1QV653TR76#V;QV2N7QFS, 
@4$+0+.%R00LQP&53&4/@1#Y?V0K-L['+IV,^!*&9I#4 
@V^4O]#'XWXW?*V&H-W=?*:9;+3!P5NW&?3_ I52N* @ 
@ZE!F,9I8:#0X7.U3Q<UJW>%%J,V%,@ R=%*/(4"C>O8 
@T8A7L[S-9-NRB7X#CO1/H?3P-3QQA\U?)M?'.4TFG[\ 
@[T- ;OM&I9"CRARX[+# .,Y"%UOWO^GFO>JJT/O73[P 
@0N.VYL6@_42WT\O)0RXP7X.8$"8H5IFN]3%@=<\",E\ 
@23@FJ938W,4XLMIZ"PVI26/4U#H "I!]WBI+L%,T"[0 
@40>RU@E>!#I#M1A4BA\&=#7VM;.B @ IU%2)U'^S\O< 
@-T+^*ULB>3\4_4)H^N7Q,5N09;*(P$=6FVU[)U)G#%X 
@"GTEZX K=%_%!;>T(IL1^-[O(!2T!@$U)9H+U:0#D , 
@O)4%14Z,<90!NBD$*""2+J0"?$E;R3R2Q!YZO:WJ:T8 
@Z)S2&G:& 5+R-["4M=A%ZT)D'2D!O\(P4KNVA2L1)DP 
@T<C7\W+SD((<RK(4WEF?+1K2M?M+VE YN6;BR?D&B'H 
@-TNW^%[VC [_H,>>KJ*>;YK0<!Z/9&%N07Z8XIQS?:( 
@;&_M.Q7.%G[9(EPN3$!^?;@C4O-:NAHP!V#%.N4T;\  
@[#[\05)/ZX%[2FU$D!9I8VT7986>Z(UBFM- 2+;,[JL 
@ZGYGM_TT_!E"W7LLO\^D<A4ZH0GP5[VFY[MLBLW]:'@ 
@N9I#Q":5L;](%2,^T@7,!./,]^'9"/.LC?[$&[^%>+H 
@;)(R-;LQL!N]LR)[ W9>,-1_TNH_I^*J]?X#:;^_1R@ 
@\_?@W=.2VXH]:QSV Z3GWZM(]13@A'=ZIHZ[0V5CCHT 
@-#[3C*O2W%*&55^G.ER!5B(#@)/'9>$*]F5%3?+)D0P 
@RTFULCS 'U*&#UG24)C.\!W#/6S7@+IX3-=]EJ2)+ H 
@2NM32:F>_+$^,^..F+TW#W'A$?D5HDKF9FV(1ZFK5J\ 
@N27-Q:%/SHZ";VSU5ZY9KPII- Z'_7%P@)N<CH*\P*8 
@-0UM]/"85@LB&[O"DC,VT!Q80<**M]>+GL6; B5S7.( 
@;-D7BH7-T9C[3/Y!SIV[4GV-^K>L(D7.H&V4?BGXF(( 
@KW[T'?6*?PJWD1D^J789<R$Y1S=/33#^ZNW@G$'_;6H 
@EAY\GI&TJ:C#JP)M\J+)>7[)\^]"L,_H"W@?;4T'DS4 
@J&NV\X_^Z+<"WF(BUF '@H"*#%A</@8&>. X3K\;HR< 
@7'*9DQ1IZ04#-SV69<:3-0H1-B6?J*K;2\!7XEX/G7, 
@2'/%*>Y)Y?I40CF.8 \P<JCVE!TUWBN)ZC*S,SYZ9HT 
@II4^&=]]PEZ5@P8$QAJ?0SBU+\A\X ;D3M/DDQ 7!9< 
@SPLR:XQ94-4T9$FWX(5BL0>,7#M-SZG S8'D^+T 69D 
@1_%M[Q]W-+'L]Y^#W/^H/I7L;($G4G_%X=54WAI>93$ 
@&BNI%EXETJP*KGU^(S4)(#$85;8XP\]C;ZYYN&(W*U  
@;N(=!"]&1&S!"<2833 14$5U+%FTC$ <J=[IB$*XM9\ 
@E<;/\U07[T[YS@N!7]IH'6[%C\&AQQE;(2X0COT]]T@ 
@&ZPFM\@/P7"FZVN(IG!%;IJ#O52V*<)D,IEAQJ40(DP 
@,2)398=\  Z&7;$K'18!-/&W1B9BU,NR# 4I/+)T)FT 
@5F(SCTE&$)"=@S,4&[GJV&KQ>!NFL(K7"B_H02SJ,S  
@5PG$=+*9*M&7@$;N(HQ F LBS,<M;*'1,9KR5>X^;$\ 
@THUQXJ *P'.2#1X7+66Y%7'R$5BS4-Y$%.+Z'QTQ!9H 
@D!LK+S_%KV$LY3C(.^12-RZYH0$Q&)5#;G<,%65/-[@ 
@O;>H#+_G$RSD6FD"4IK5&AQ_2AH5J+0&,DX(#N_(9N4 
@=G"\VAMG8N3E.Q0B3 ZUDP)QCK9CR.JQ)9=R_WOTEM  
@HMY-^FS &L*C)M'H93R': 4:[0?%I*^<ZTJ&V&TSAE( 
@9_)O?]!2:L3><<.9L R N52>$5%(KZ:KC(DQ/O">M54 
@7RZA4W;R@VSN/TSV*J$49(/=UEJ/JMA. ,<3/AJ6YQ  
@42@CY5,JN7%- 0'6UV>!?.3_-!V,8=)VY)Q"9^7M'<T 
@E).$N:$Q/HHMQ7^MU54:S>)ZS# %"\ 1"'U[=W:SF8  
@_TK)EL:&=0+,(7]-G?J-="MI2.]7U5#*+5'K'E9!2@D 
@'$7Y#WD=UX^>J^U7C*NRV$1,HCF<BIJ?\]_-!H_^AM$ 
@<\)<1 ]5F#7Z;]A%(BK4\.C%Y!?Y.M5W]MW'*AN7C"D 
@$0@<G<_)TKOC?MHT*?^,4W75@PZ[I$8EE5SMKTM+96@ 
@'QV](^X*X^?* X5_MK13Z<'KOV&[Y\X&+4,TP !)40  
@Y)IK?MO:*?G%G*P!77,!L##$4[$_WQ,CBZL"O*QC42@ 
@<WFKA$&'OG1EZ'Q;OI72MFPNRPE(5C_: ?)YT;.8MY, 
@4"_1CL[(1/:9[M?O>?+;JJB;>\0<=K2V9[:!G=1R4"( 
@866"C<A>CBLM^I>?\3Z45#G-.$#4E_[5@4S9GJ-H5@X 
@"<#X#VSV3!FOG49R/R-0]G1JCZ6VZ)M;R>XI?G&[];T 
@M4"_3\KMOZ# \\.((S;Z:&#&>;,N5CL1[;B, *X4]0( 
@/N.]L/<<;>:O<9;9+94W.:W8NYEPJ!,PL6P_EQ.>&;@ 
@V 880:'"72<=O]VQ@JFTTQN/F8#A;P&9 (J.&NEW>3( 
@(,_S(B$C1@B#H4AXDW&7?Z!$?X3JC0_='T[81^[L+S  
@0/V>&EIC.A@@7^JWGG$8TIH!.#SMSB!J7^G'3WD)SLT 
@77)Z(73?G\X3D8$<  ;#,Z?#3Z;4LK]_17"Y5?P!& T 
@#PWE.-,D_2N!3L&BL/.,WQ%9*>R <;66UB].X+\[,*  
@Q+KA?C?JACL9BH/+\&+@-C2&!,MBQF]BUE_8T.,E1/H 
@_*\3_=EN"0QU'@1/'RYRBCF+6J:WE1OVZFV&_<$T4FL 
@0:[;2C0"^>.H>//5,M8^/\@("0F*XEH9!H[X::7F&[L 
@&ZF?(M<)\6^,3C)KX58OW-=FBTY/L8@DOMA.W[*V7_( 
@K=G.[;DJB^78:MZS+4QFS88T"Y#P+YOJD"17U:Y@N80 
@?MLU'<%;#!D@VKE;  @2/9;UFB9%>(7=VB@1VO[WUK( 
@Z'T(7Y[-18QV(-?XD>7VO/!@*[XH<4\>!.;[JR(B/8, 
@3Q]/"XDW)K0/=RBZ9#PRU-0<^4,1.3!Q4=+1>NA?PO8 
@@CZ+Q:Z/]R_@WL'X/0$+N?!8>/\\/F\)%F__V18EAP  
@U/O,1 ,-^>TDW)NGIPBNOYO1U!Y3[4C$'+7J_?RM%_H 
@LQ'.E=+5;A;!1X:L(I'&+F)([+,CS1E*_-!44#)<3%\ 
@O<8+1SGUF"7X=?C)D]),H@Q2<U&X)B?6K)2)1=6GOSX 
@(<;DX=M?9ITVRQ\Q5ZA)PHPS"A]T*]BK5I16$AQY(3H 
@"$T^"D(FGND-78O)33<F!3A_=\45>[\SS'\4((N8_;  
@"=C\AHV3;<TCDXFD$*,Q=AMX<YWG\XMQ'[<HOR5+A<< 
@-FR46P>53U5>)*8IT_%'_K183YLL)2QN1N?HO[2((,@ 
@9*NX""-YQ*U>O11,MC$Y)T4M34EP'D1@1A"'Z+WH,4\ 
@-AV+T% *GCOJ[):N 2[HKEQW V*NYJ\ =WP\-U@?*>P 
@EUFL&(!J .&5#GDKTOGF21Q9>V=[OIGXW/ORZ5/$@L@ 
@H'009O9&EM]?)XT_+%&%3I;IOOP-\[,=Z*]0 =]+:J@ 
@5%G'"T?;.]Z7;T;:C$%;=DJ.:$OS8^^;,%<!OE_;\&H 
@3V>+7-SU5;""V_QT-<(S$JX=<*&']CA S17RY.#92&( 
@!23R*4#LA[3C_D'*:\;T^8WF\*(&#>[-C&(/LAHDF6( 
@K\;J]>I-(QO-RB;&D,!V3J-6O_5!,GH@RG=BMH7$-V@ 
@^4U&WG+ 89S \@HQ#AADLIZU,*0$W+'_:AK7MS[KR20 
@HO!46@[EB:].7,[WIS@DN396=WQ5K&R-VZDR;]^4TLD 
@XWJYKM3<*,=;VCPG?Z<]"%SI2?S.X:9*Z$T1OB:G?/8 
@/T8M9G7$M'@I1P9^KL]47/._?71OT8X)T%:4=->00Z$ 
@4*'QY:)>EF+JU]2S#<2R<RX:LQ^0WYOU@EB-BOYR\R$ 
@_N@?A8CQX[S<KZ1I*)-ETL;ACLKV=*Y&9,=]0S7_\H\ 
@D3$%51JEXR;=P^9R^<X\C6OHH[7GFT(XDAIX;?G4: \ 
@EQHL2PX.95'(=NFO9B%/'>R(!I%GN56/6.PDIJ(3:KT 
@5^\-YB<Y_^J=K-Z1Z6SP5=L4H[0-J\<!"A;-X3UZX[\ 
@5??2P'^C=&80J=3]B-*XU4:A'&^[(^Y+!6 9L017'H@ 
@9FO[XT$E]W:E ^P@4R+J7?:?8H%OQQ6YE+?PFH]9_00 
@Z))2V@L+QNVMM0PC+LL(EC4 MM.<,[/O5;R$D7;W(EL 
@R["/B=X7[S.J4Y:H/71NXJ<A8MU@\*('6\C5=.WB 88 
@VD#E\>V-$=]1YZ!7\P\&A_2HN4[L!V8!<2KZI72*G#$ 
@ <M'@ A*ZX-$(#D*?^L=F>('%U=BL'/6,7I=;'++5C0 
@EV@$GKK;ISEJIKG:\HJP[?[9)P5ZV;WVYEP@[%1KU;  
@7AHNPDGM]E]_.S+;Z$(T>02U4(A8Y6WYT!LQ_! V*M@ 
@!,T:OPKY+4J4"C%WHWP.U"O?!/#LVQ4>F[N#++Q:&]T 
@1^$WI%]HA8*;YQF"L)1USNI7&^+&P87-::P@[$H7Z+T 
@[,R4"82B3H.UB(G&L1[^V;#3KTUF53DX(E[(3Y(IUH  
@H JVBX,%+N;;^DIH(WPZ97J_B[L<J>JIAE'VUFM*WS@ 
@7,CB=F#V+Z<:XG:SCXI,2;9[),# JT$GOZZ)"Z9#?U< 
@74^H9JWSD+9]XGN").1NYWZ0R>C0+-]>?4("JP+)JS, 
0G+7PN;[JP0%VMA9+YI:HP@  
`pragma protect end_protected
