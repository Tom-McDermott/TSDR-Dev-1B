// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 01:23:35 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qUNhcICsROgPOOeGCPl6M+urpSZuqW1wKnKR1s1Z1zVaEL6fkML4Wy+3JfGfvD3P
tvGdg3qwT7ZCYUt5+m26LVVuwQVkqvppfV7qXuOoaYMb5poo/rOPHMrC8xOKLaI2
ki8RAZs0fetGABjtwHiWyPQyus8hKSGjEZN92kYPPJQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12336)
FFafNYaDfKlvFGrdUBUEW3i73sPcTqJxHcBwdonFS/VXzQNQtFAm4qx18K4raDWl
0VGxTv2T2kOdvC/SqWTKIvcBaMUyX29R//bPwVT/rynabomhy0JFG2kx8CCR1tw7
46rN31cMlAkY7BMkndz/COtX3R8F7TxthruSkHgDl/W6eOWsSGLKwoV5SfYK6PjX
Y4RnNwsZKs/tZy/3RljLPZoBSY/Fy1WQCr9ZzEzFMZUFnvldWXoGi8TqLPt8TkBE
djScq0AN0RInhIXPDMCETvuqU51GTRBycZVuhFzJIT1DKiXiDkiBSnsZ/s3WXDh5
kqDA0k/HPXYgIeESqo/Ypmxav9ms1n5fnS0zhnotzgpd20QlWGz/+L/+nFWsodNw
OfeKB80i/QcmfZgj1LfBLSu/ojAk1eievINPah4nJvJAqmgiSiKWAyNka+yHz9O1
0X5Qcxl0qvHheDWP8hXV+2nsGYnS6F7op0qJhezb2FPEhevhyzvNwEXQI1PXMcPx
m9x4uCvOMZ5G7YnUUQWVu/AfebiLDrhYr0FwAGX10q4IjFjDVfFmDcn+F8Pi9DL/
ymi9+AIYImp3MwVODq5jaoubWgL59vD1+dNot274FtSaX0+1+F3Jk7b39Z5/qI+L
3fsI9sx9JdAwGK7J1jqBORH7aieo1o4YcHhv37USNsMEx6VfvkdKEvrveIpJYyYi
uc3PAHho9pAvqY3/pEUofwrz/+WFjUcZqcmcsXRcycU2kyvAp1NjZafwgllBcl8S
vwNRAYn5u1PA/Od4DVBtKSYRSnUfW8KRQluybKjlY9NMKxlz3VyFJ+iNHepj6h1D
a6b+lnDdccgxC7JFNUkbNFS050fUi2iWGNQrex9evmqZyCoYQsxKOaOzM6O2Wz09
KuY7lGw65WFgeDdkd5IMosYCCQuJzAA0Blk930Excyt48os8/7xzeC1b2DHtq0kP
uoLxXid92r32nAPSjm6Fm/6VjvfXZoGe5aF7/EJCN2eHgn2kJG30r2iR6kofGSqk
gTON+Qc9Tz67gfA5qp630DN4Uhf+ABc7GaX3yfURIuUdR8mNKWWFDlyyO/eNulG8
2K7A0shGOwQMOFTmI73Pld3oiPzFRKUceR1lsk5sWG9vDdgiYRLl9BaGwl0i/L+t
gucL1YFGGYkZ2qAVjC29fmD0FFBAiVy0Ci5jW+h+Ml5nk5eYZTNWxpspZVapnwPO
qgxyKpczYN5q/zvMixrcJs49fPmxXdWQ17FVl/So2GkVFNAVZkYE3RHp6Q3DVvwJ
pLLZt2sc+JGWMy89wKHeABRx/XB9i+fIXk5yd/1y8x1JvOV/QwYJqaKO+LeefTje
Yhf6nbuxNml0pidfb0M/LJQ1p6Roh3/GLopWZ7VdYqMP+hwASlWkxQKEDl2CD9W0
+4QM8ixhsjtvQ4yCqfm50ZLaukBYOyanm0b8IaOtLFNe9HdnZzP0dQyUUavCZ4bU
gDZeG//Wrlbw7tf/cqNj7CzaBqc9eI2TMFesrUSiwSVDq1FIY6TAqxYTsMcuUuw9
8Pi8vJFqmITKe/KAUfUf5T6133Nmld3QRyL9PYy69QDHROGg0FQDee08PIOLAlzE
Tjsxu9NlUIHbJkrI68RnwClTrRe6WbYljjDaVrvxXMhvKary2hrA4BHMll9UztZc
xi/gtslgGEu52sxmGgay0+E7lNJ6/PG5lTV7V2BwOoJLlPWLno8W7EKJ/uTUb/fI
fAaMxoT+0G2SqfVta+Qer9IZIrWJRoF6PH2B1CsjODK+XNwaSWdu8nst8XcgA1sr
E3MiVTrXBIeQURlqbm46X8D4uGuBBZXNDtugtYUxhOSu0Sv6t9cvQto0HZJjUMvB
NHWAg8M27OpHU2M6d5Im1pMYHuqaBQuxRq1xADPkFmmKaiCoPBU4GLvvxpRjDEox
kQw8WwVn0XVlDWSIozvNq1Gl1M0eO0YDoUqIlf1JaiaKcBumAazqhEHsF+aThVVf
k1obORpreDdqc1kgF5axICx2JsV/YozGC+mdyaTDvEECxOK6XZtcoa1jFNeQ+HWJ
ILY24dUj+OQmjvh6xdIidwFbOMFNxToNgZqct16JAMkyP1ij7muFiikxEJ8w5jOk
5oxHP1MCBm0nThCCMlCUdZDU62/JZDyB4wASnvhb0MI4233giZ7bktL+8TQbr2LL
pQvm8MOT6WRP6P8TqoJaGJdzbehRfAKUA4q9iCilgO4qybEZflkOO+xSaphJyEzO
4IJkbBb0QwhWizHSNa/2MgIJLCLZHagZ+wW0BkjJCnIEpxkDQ1Sv787fpXC5kV56
qRdmEaFmWSxXoa+Ls3yeQ2ioR1onwR6HBWfafAWgjeFtOgiL29a7V5SJ4Jss3/60
jWm5IJpHLrPzaDBVOrlUgvHijUdTtOn5zyFpInHyfvkXqASJItBgyAdy96BWIBuT
xEH9JNMuhsectK9d+lgi6JDtFASBaxnJkfMAaqQzUsCZr+zO9ZPcmtLNF+/zlQOY
OGT2LuwSdzW+84V6PPFHtsz5aprDZhxL3yOnarvXMfqYJkGaBYZ6hkK0ImYwlzaM
+JWKpq45BwWqOhzpMsSzITfn9SG0JHIfTBupKPICjA+AdESoKTFO7StyExBQAmsO
J1B7oH7O0DcdQsOFnUsSDnN7YZvF+6B9ZbKSOLr+xy3X67AzNfJN1breej98todU
cxjymHH4dtX/6Gw0TqNdtxubjga+tvhu574RpOfX1njOvUQotDmn8cCHGzQGcvz9
eLw/KkrnzoyK82YHfVQO5q/cBqwMAvg8UNWcJ0a5os2ZgBr2mNkpBExb6JOhuuYe
L1vROp/DFjpLurNGrJaEaDu1X5SZhpUBRkR1ZaZHSLtHNcxHe9AeCU7aeErS+rcA
6CyqQOLv2GCLQ3P1CS08Dd7gHgPTzioDeZTMQr20HfYdTMLrmrbj/sZ4A9SaOEj0
z/hNUPDIMTXNN0MOdzmfyy6e512lrVtHh3UcjPUo/m+vjSnwqMlXj2NIQmsgizA5
gG5tIMCfrccWOfy92JFMqK4Ta8wpW3bZiFJ2IsY4qFZvoo45psqu8HQSp4uhGp7d
zCe8YdJu3b1BUWpq9MoEPE6f/o3DV6tEWtH6Of+teaSUP55C/J8yYzvX3rlMZXOB
iGRK5DNNLRigGncjWlCPhPL7WIOuzem12+qbeQ4CPRv0yQGyW/N4irWDJE/p+gr1
2QPlAnVQwhzmQt/l7801KyGAUBgDleeFmd2ZUFqGglu6As0GXhrDbpW995ILQtW4
e4ECpKX3RVMZNTZ3EaRik3YkVOy7uHRxYHq3YQ+MeGaJUpuGSamytinupaFnOig6
0o8i4mEWSFR/I5d/I6WWNbqvv7mtcYhmUwt4t3Uz+HExAV7kitCuXqVB9AQkprnX
EN6MV50BslLY46+iRRuDRlI25HGK8ysb16cJRCfWIUjdQiqCtKE7Fkr/5k8ArF/5
A1E9FAHom+byYsilrXshp5Sma+10SuL1snFHaxqiip6lrBnv4Tbl3aZ5N0+vavnD
R/ltgwzJPFfdGCZQBRLsH/GdWyo2ylDwUe4Chtwu/akNsu6piW8ujIV4+d8frMrd
myh66XNB9GJtbouCvVM1c8NZxii3vxY/OMD4C7o8X/VwIOP2u7oT72wOZxhGbxL9
MqR128hArnLTLG0BAp7EL3CocNSw3NdoLhuChy0N+z0mlfqhET49s8UwVGS2OZ/U
tV0qn/UbiTKCvOSJMYcViJx7y+iYsZK0n3YsBerpSfIOVhzPsBNz4IEGkW67V7DF
UJ4PzImpol7M7vLF59YbcaYbTZAY1/9ZLeSAmnoxlOvQabIsUH8hzW17qKYim5IO
h4mAOgw4/rqvFpW1bp6bzeZlHgBPaYya/KJkBXyM6EGE1qaUPSex81Z2QqBq+69I
ZAJsHPqajgVlE9dO+ZaO2MobLsWrFq+RV1OH9xtoHG4pnWQcHJz0iEYuFU05xMSY
3hJn2ZgviNn4EiygcaitBmnZem7uMRHeSaCPXS+1wGxEW7oZNyxvN/uAhCJ0fcu2
YWm6BeYC4jB/BNoyJoDhq9hKWE5ZPHXHywM1maJyi4QfFkoPNLDsrWOPlkzkxViv
fVDSxst2gRwcAlpbTg6Fl5iDlBYj1uAIUs1Zht/15xR/GR87UJiDXBYu3poKKyR2
V/wGjdC3Kv1vUwRKREo6QsMxr8xQYtS7qv5r9WU3gzjlN46DhEF6/jntIlhfy/bn
b/0QjTKVW5dL0wb1cUHVAbYCr8G/lIu4UKdx179Q5jlM9eQFcyQta1Mpsrk5smAT
ypNxar6sEDE1xq8za7hQqymvG7eCFu1xJ3MLCX0PUk0m+Nje2mtTgc4rDKklBxT/
vHQB3FpFQdyIVuJQJ9lhMrEjKq6TENlOShPJYAw36HLXgtdwtzn7jnlSdL+e2GRr
SzG63lDukKTlDKMKRFlo93FA/qq4f7+SsyZj3z10rBYVbU+wwPfdOfB9oh6twHIm
0VNtMzW1SxyA2BIevCipyDumUh56saNNlFLXydXWF12aSyZzt68gkdskKCnsY0KG
4wLhSVEiVj8XtZHICG0GmG6IKkDXDsCZ+OP13GH8uVV+Mh0gGbv2JcQO/QpH3MOr
hGEwl3bQesEM374U8o+qapgN1m84KcpK/Yx6qUhdQ4X3O2sTLWPwgQ7Tf8T1Rg8r
95DNoXKbPsr7w3CNm62zz0nAauXUDjnb2KJBRWENRmk79tb9ZTUn2c4I3I4y1WaF
B01QeLkqCoZjgZZpWMw/4VmDrUzqzPivqqQngbo4CIIT0zzstfXWF1enaBOmkY0G
vsIKw+8imcuu+NZp7PtN01Ci3zXc6dhvAI1YEWn2MuL0ytTapZ6hqJuueVpR3W7j
u0c4NbC45Q4c8bS8w8hbm28LAq4SaTcA+KLSpmMnV6GKh5Uyk0wsEoE/efZN/yJM
UIi+g4JgxragH/HtVAzrce256q6yNs1xpDeFSz7k/ee8Ox1NCFkx5Ze4S729G2ip
3QaAlQPcerU8FYIcj3356h9675sVDDTrV9zKZTgh/d5f2ie9Q7mU1dfg3OAXJjQM
ewglG5+PWt0r2nLxc0DGLgfGnCKxi/hS9xulQQq7g9ajAdUYK75JYZ4LJxGBDWgV
wYUxwaHiiG/7lyV1TohWbx2bFQVs/69Mu27Ct2IOlV8g3Ht8t9gO2APIZVvUtwS6
pmapatuHvjup3xy/wqZY6G/nCzvGJaXCl2s5nyigfrRMoShXoPQ7uTT/QnSFJ95B
mR0OxilPcWVXGXEQLkcdFDVs5xXxijuLQSmM5uAqqg8uouiaYIUDqS8fYkZUJt/u
Rgsdi+tdu4kelWpYthoB9DVLLXSNAtGFQj/lp3TySJhQG0ddoKFgXgvDcvlBwWNF
w1lJbICd9XEIpue+BPz/o0eETMWpM+h9xCsW3i8yZ/2xq6d5D5lqxS90GqMtRsr4
eGTRzH3sz/92oUmOG4WL3xEbCCtxwzd8rYE0GMrhZtcHVoZ+9zhHB8LwKwS/+tb4
306N9M11iMRrkmRYSDbX2UC+w9Zgu0Gla88KnY6sSjZNBzbNcTQRnhBlcVxYnbnM
+uZ1gNsCwqH64TbTzzWuW83W6T7Ss2IIqhD851a55HY47inloGoUlvIeTqSLD0BK
hYHnpnF0ndr6MPlMGVshaeoxbMZHeaczzfT4DwSrseNbbSDvSZlV7mcfBpJYzvSC
Y2cWsxgtMQbUg3HXJOlaUNterYX+F2H9KNNfg7hTtp8HgE73dMwT0uYNlxEP6l0x
P98ZgxldTVf6ynB7NFyKqiHsZZf0IqZ5041m5xjhCWGFUPVVZ80yyFpQohKSCn3G
rSF7tnTjkkXyMPdRTMm9Z4GhjpLpuS4tdCSEOR3ylst1j1aZmQAk1lZeO2nPsVxk
ys2cFNu5OGzJuK08CCMBZ3wR/Yxce1nNXanzv+ESczGglYJ6qZu9DcYahdKVBCvS
dE67KqyIj+exyAAkgk63ZsQkpREihZBornzdX26FtzJjB4F0ddskhh58poZ6eGd4
TWa+lT+8zrsOAvLXypV/r8WKKTPtEHN5EQ2PKEjtOFClT1aOsWIdGqREbbNgV7LN
sqYveNfnE7PGOYEPZppKBaii0frSbBMc6VdjBMJMx2DqDvxDEVsb3aBzNj6Y7Z4v
VhnClySard1wnGSBotcqmsFjcR0py7Y9dSURJW/Nd5S++xEPDvaHnK3aurHVkgyQ
V02mKntJw3AedlpVbLJCTNKET8rYZaBrOCXjDR0q8s9PaAyISuHNff4AHDRoycRQ
nEHz9YWLADrMlq1teH/GvfnqIpEgu/98ZHDIMkdIy5QEmUZtT7Pm8jEP2stZEEw6
ykvusckDzPeBEXqS63LaGUuriTJKFOubd+lUX+sFnM31JvkPBmIh0405+e26KAmK
g3kCriTM4C4Kn9qEqshmK+Inhq8zEbtzlkhMoOohRNGD4Fl4GFOncYkt6HVuTjNr
mm5Y+s7kDWbrZjJ2cSdv0VVq6yzxhPMDH9bTK+2u2Sv/GCHpsqL2w+a+bIwsbRd4
FYORwKlAu0bVVRWgvlZNjGA/qpeiCQCPzIJ87rfEcKmK0MubQaUjBMhYWks9Z+DG
9e4oJIzh7aQTY7gGOpADhph5mXcQdEWPMZa8sN/FDaW79o6TpmPbtiSWUY+dxQc/
NKAz7mED3UoEyli7YjmVkygpV5o4TEL+IG1Fd5hR3vpbX2taKsfrQIuV7nU9g0z2
pfNxWipsM0q8w/lbTs3Ppb+n7u/1NfDK0VtotIruUptvAg1woh2cyZn82SLKrZzR
nUXlussBJ0y/TnPGUiP+6UCVYnjapn2A10WXQdAhuW1NiMxFcrXK3JKBn4zNdUWy
W+RsC27Y0spCKj4gsO3BTGxTCqr3GfKEYJzmUqTzGgxIsgCXdr+uij4lqPZBEf3x
4oZicauYnihoE62o+6nUY9H8nwTBR9txEthDEE6fbIbDtkegKjFjCNO8J7lbU8JA
OImyCfs3NVyCagZhMZCkMR3KYXaPOeT0wHL6mVjBFNjp2tgO5W4t3abUjC9I7VXa
xKMMLAyAfYynTI+m7AsGPU/vFfU7oFRwd8isQMDFJ+q2q4aqScgndE+FcwCzehdq
ws03uHgIR6LJl9CujSY7oBmIyzjmCVBuD8Hlkouk3PivCdX6O4LYDZnmE75e/a3R
oc21SBjP1a0MFKyf56/amJW200elxTIJ22ubjwy0nu/ZNz1hpO6zpWdwVYLjDCyu
hDj5hVvb9RM8sy3cKo5tNuWmoPvq+52uy4AObjEYjQqE51xNbDjREv5Z9wIU7q1M
q9TuKPK4OyRNmtx4gwXOrdYr1NMp8YWiIlHb2cHDn7fFx5leQ42kJ4agS4AFT94a
lSKTJ1fjqI/0nOQY6npRvCIurRuSKEE9B5NqkzSW4v26locLG+JrQGbx4uQx+llY
7ewenCyCDfPdi5ZE1LAZvf1K8t9hLB8ANge+bQzpNkmUwma6nz8Z/ITgcSA7JRUs
ytOCApv4fWTn+z6bCo2RzAM2AybwO8vpMUUfX5f+p9ZN9h3waVrFAdRTkD2lWBZL
JtU4bllSCgPy04BWQ2M0mO8291BpxCdot8VKozeV4k4QTOhlMyyhrSQbeC97llpX
D/JsN5vtux5wJN55rn2Js5mCAXmBpeeLI3qOWByD3LgAhND9+TUfo4n74ddVOxVQ
YMGYAcGyXjihoJSlEhDPpK3HU/M72No4GMJyusyuHqo2N3KrvJqtUUctnf4yn8mA
/G5sYIALj9FOK6QJVsSRNYVMguRJrVX9NobTyaavsKd1HIIddzJqWJgYzLxHnHP/
rirMv6OT2CCEuR6sJtLVeiIV4zqM8Hl5tXjdcNW64Wp5sHoEPwApIG9StK2K7jgy
esY/a2MCaC9EbnGWHNWPabI9XHzucZcvegzPylL0yfDX0CDcvIP5X7tkhiMmsLly
1h+DpYXkOrOhu72paziz74E7kehtRZiBqtuP4yY71Hw9TAVlfuyrsPe6kqX4sXE/
O5KSWM+HOI+zda0dqeeeNU16zsJp7HDKXV93dwrXh58KR6TJQ78mt5aqcl0Eoijd
K1H98YP6ioG4+Ln2Hv3x7VB1joir9nlpBUwbAzBIc7H7tl5Cr/mlNm0X1ZFwzglJ
S2n8G9E5yabTY2zWDWM1E5tIhTbXtCOIaB45aTMTBC7k/bQdg0gO27nAwE8l/4H7
HAbwayE1Gu5LATmnQD/S/c/qto01jkqS63GuaYrRCOpxLmunNpTS2gZdRZ70isPa
EWZRbcMxt/L0v0pxZ5sMN22KrhK6Kc7E4vN/TOP2QXEVp+jPNIifwZNe1kDtiMvD
FYN1VbIDCCx5IHGA2KTxSTwJ2Yimc53uun7JvbKvjnWgN+TEAH1tPxzcS2lbnEF0
RQpYhA2ZPXzh0NU5zEQVPyZC2fL6nhTkrJB7xYh4gcYOHTjuBSpwKA6H6USNaU67
PEVeDtDUQ4MDatH4xVSx4ThMglZwheoODJ9d21n+MuC4XhRomDebc2EOLg2GBfkZ
XO6CuBeYM3XGAauqbYlkV3oRYRmq4L83ZqmL8t3PNJW4G5GQUlSFdVV5FCIbXPiq
O/GLDthxqul9GOiDQPLk3XfDszOYkZQZRvnn5ZQbzqihWjvnPoW48UK4zdFzPtU3
BtA5xk0iZDnxjngmi6OCWvTYjYxFqZa9vqxBX2uXqnCsAtBsV0dqlWmL/hqtrrnv
gDl2z80j/E40m9vta9v2ad4RXANohK4pWU9TeB2qd+vpD+C9rneKWeFFMBqRe/lV
dXNXosu79TBinyP1k58YdyT16ADXgnLMa/lRHSE7W4vHdQJ+GhBbbzlcESrTmxkW
MqRu2QWJLDmRaRgjihxU/kxIVkhHolK3+Zj7VMjJUG9+EMooiSgmRloeDzr7FajY
D7qANGWL5vjAzsHDyypDGAyZUvdWHuP1xb7fbGo9s6NNclz71tWTrKKbmREDYImY
bY1RgGzbCobSwXFUUnJJ7N36OwuEw37XWDpVqTHgwficCacGV5IWmNrNYSESFi1O
saYOpQU48/k4Nkf/kejDfi1NIF8qL9WYxeoGcODmLfe40AzjtqDdY13FoB2Nv+j9
jA+gP2qZ5VxQMaiiEnXy6bkYlOHr48oLrzoWP2Hlw0qbw1S3E2YoulI5ov0XcJqq
A/eRVPW6X6w+f8DH09vB5CQba59kmy+KX8tnrmbhJHy3rThri66XTrFMRmm7f2WF
dwH2+Rk+faVqgD5juaOHwwphajBtn+v9dhwwQDET8DwGAwTbQIP/gzQJLek1EoGa
jssnEu4L1bD1jqv5XRE7Zaev5jyZEcN4rRZ9qEPuvsOUeQW4Xnxi1HXUbQa5F4xt
hrp2rWnKR6uDpK8hyDG43Sar8xAAcyCg2A/kKh9ADUWoMGNGyCEkNfbHErvUWvxq
nptL41nkwL0m1LP8QBKrFvmf3cRA+Ed4l0wZe66Ze+Ezytbujy330I8u4TtvbtQo
LoTlTjZ+mmrbC6i64GP4I4VDx4dTOWGqAw/HS449hI0PwLzJJeAepD+wGNrsDc9R
V8XFNGKVfoLhcvVbEJs60NNefPahKkEp8hVZ5Xj6EAlMJSjiwlufNtKgBf/2bi2N
Pe7q7stZXyI/SVz76AYGWnJoCa7LCBiwKOD1hnUIFOXCrB7aLYmdxXQPn9oVH4rR
2PUFHKbu7BAg1Am3HpPpC35s/jf8uaAp+vnLmcN5B8epZZWoV56KpXGmudJgOweX
MV/LcSKlgpuC4hyx3VP3PSHrxUlInvX45jenlhUsEnUBLIwzd05MNNe+6E9NSgrN
ycQz2mFMjW5w5infbV1ej+xBscf8pxxbv3s930J11jQEFI1wDtJ3RW9ukKSYCKIR
TKGHxaQVnkkPsMiABV52xf/f8qVsSuqUx/Oh87PRGLbuQl1KSEaUqQ/0rPeLA7YI
ywowB8bAn44MJWTMy04V5dQWVhMyHtGC4WpMltJGEVqeyxGtcDfZUw+/fOrf04eR
xCzp5G1Tw1IKbnO4WWlL0HxPPicN2gwZGR6iLbC9I5KaKbk0tA26kfqHPehd2yXM
dg+lHA0e4GDEvzNL3O6j7F9A6+RZhlcNs7nOEiwtltk0ZNpsQal/ESDXC2FVDXnz
RLZYe4LdJsrZ1xDyBR4DM7GkOJkY3LC0wAI0r8dT0A4tjMIVsmSb/inR+7b5Zfik
spnD0FW7eEDNWREd1U7u+n6LzBhvSyHZz9FmawOMy9AFdWjEpe6xe79v15oPWpsH
o7RitCXSBRSUgyTtkIC1/H5tD2bumnu7jar7bJX089WEyvUKr1LsXorMixGXkU9d
Sd06EIhHliddPVTTJhuMZHcQ1+Cfk+hRplFZt9oneLLq0/vbs7kV4N2OFGOPGGIL
qMyzQWT4pVgBZ1uGcPIoUabyVESsndPyKurTL8lg71Jmt7wpRClBHMp7JE0gl2Iu
oGdy4N1IUfI6PfAxuQyxb9gYvVs6Y+vgG2FT184uZoWWH9b0UqAc+oKQ27BDGas6
jpFlSW/0P8y4rBlfn8sIDtPnq1K4yZ2QXuG4VvXZ2WIJgcmZyWvEqE4Gf0X/XbBx
3N90qaFpBxU2tiAiF3pKzCmeKWM1G01UXPmFQtmtjd1ODlyC5nkz8+MCoTzN8+TJ
41VnlbyUnhamuQFkH/fGhmaT3BmGX5N3f7deWSinHGZQ8VwUnDgE8bBTPkCiCnhF
BOFhzzm9I5NT32H24+JRaIbezGbkuA5JGpiIKc+GVtN+0zAKwLI0stC5RqEaQM9S
BB9YvB7JWj2zzR446fj2RARHY0ax+wFY8VeBJr4SBoPBvkikkILa4tHL+tqAl1h4
Jnd+u3ErFro3mb5qvua35thlursgbci8rfqheUm76eYurqSqC2TkCRorCM/ylelg
PgDbD09el1Wf7lubqB31e5gxSX9lOMwt4cO3MQLbrCYSj8hd2cIiDejh5K0V7is9
z2XF/tM3Ko5Qo7LegCLsNqmIKK8Gos8BqI2B/n287dAOMWOKj67OLdIullxnyBJl
c/RnzWXaT2IaWk4v1m96C/77N5JPCCkxsL+lOHtbe8JeMiVUggyKFxSpfH17l2VR
3lSkkXiwcBP0kXUiJNde76rAO5CCH+7UL0C0p9DYUJqSchdKrFxL5mLO2HfBuCd/
siliZ0BoXdFiM9xTsL4MRhVy+kj8KsDKZylbaZjitYEkKG6fGU7fCJciwwr0wSLE
keU0iLMifM6yi/+S71iIgulZ47i2mQ0nVyC9h3jipPVG5zr2DTs3VwMQrjR48kMK
cocuCh/tHMgsrFTYR/s/0VxZPe4Pt5hSCPcUUsuu++X6MCuwY7Wbz9L2XwBxjfDc
esvO3NEJm/L9tCmjEQECbopO6zE8Cknd6TagXvlPWLxLf+oOpPAs70Nx0iQXSyPy
bmnvHYaFmun8JiW/LLhFWMpzv2ShF10ctJnwkZjJ8lvkr3bCASPB13CoA96y03VS
7Gc34Ays9nZwxn1u6HMzFF4oCQLOhmrgcFiTCgGB54jZRdVu8NT27lSL9m1uJlh+
akVD2P+hdNFYuAkfwKESmX/G+Evq/DpjpFmp2c+DLcqwChh0gouTk5dXF16mOHl+
LFqHj9PIgK3OPKJfRQISl11GvHMqvpqOwjbjWwtuIdQaFvRdkxTZkrWynQ8DlNPS
qdO8rDCWHlXJAgybGMT+3mGNmYHsBpcCSEjUcYfhInNQ+xFXkLADVlPB9D57B1fz
EpYCpC1ZY5XStvvz2KPWWlBWExX2e1mzlHfJyBma99zzwn3OO2Js/roe3JC1BY1v
J139zBek87Js6Id7ofuH+FuPV3FCyqwZAYCLAA6HAIb3GWeehiZpkwu9D5MBFtzA
3PPKTFA31jj8gqCcvH02CNQx1Kyxl3MIt1pE0VuZqqN0peS0wu0saEZF7uH9xcLr
fZ4YtIH0cwqFYDb7HzE9BL2IL08uhB8iiLKGX9Eqk+hDahKk8+HTA34hDMNVYZEZ
DdL1mCZqG67BxItftALwORL/OUMgm/cEPXJcBS6XthVft+6Fc6TWb8+L8qyOj6fq
/N0r7zgi6G4TUTVI/OkBHP+kRDzw4JXTp4PzEctc0ZYvU4RfNh5OOYhrU/FTZUzn
mZ6dc4INfCriFiAnl/Y80dGOOOcA/U25Y+L7FKNX70F+Cog7XgyQMMMmF6FhLiH8
XLlg7BNV2kT6nWSGh/SeRlkUCaAD4gHlR1qzQwltHfUzoVYvUfaUGWjTi/Dll7bJ
1HUwOH56vfQMYXj1mvgtdxz2XrSQi6qDk6s0tWyvFiVLrqD2BnpKPGOKloI1tPNA
u7281P1YQXz4cXmFOGLkvE9igSwj7PfLoSfDrxfnNr0x+6o7Mjh8/vquKgoCqD4E
Ti04gsC5cJzh5WkvuRn3fM/Y9sErw02w5+96OgzXpugyH3/lh8nDWXLVb6aowNUP
O+6v+6XGJC+RskeE47KDnGTQBzcBuwXBKVQmBSiCAT3/lNytVcwKo+wDooVYgOIT
oeo3re1j1YK3/bmXhVgClO76z8ObQxBiItPl93j0qgKivnayGsyX0CkH/+cd/xqL
SjBnbtz+2C/MaUd4U5EworRotd4ZxG7adjS7f5VXdzOD1WP6Jf5sXWxkYs1/Y9Pb
cQ9+dHoVKKOehlxkf5Oa/IX7CbGUeOXATJ02lh89mMH6/1tVberhPzg3kLbiCd1z
fN59hSlBIPSVwfSgrrOgXH7lef627fIjAftZIpd1u3wrRnlF/AFftYekR6rv8XgS
MCbVa1iCm2VvwmB7M20kAHXFDTE6VB1DdH5R+oCdNb1dCozyA7Vd1Yl95NgG3+fW
860XqTGz0EZAWSEn9AG7nEYHv8jeZ1QvhqgWe33+gDk3C5F+nO0ztdYkOaWk87c8
KAndekRvcoGTF8TeOaik90A3OSDIzGriT2UdzlLvM72gY3VYy0R+VZbS+1aSwCRl
irzJowJssRZ0pcUJfkzkrVOvqQM/KcoJB5CwlDVh5lXnJbyp/TB7BDAzNaFczXr2
stutKCswgDriB4p2d3KkMdIhUZu/dAk4mrdDFToFGn7o8+2z0/j3NvZXrbXM4C8O
Gv7maQcjmf8SNSj2or3L21cN6j/bgtyTedrUh3c+I5v+DN8+7UgnmrbCCVNA3GdI
2f42xDmGv/GIDrfU+B0s8E8CUU2EJJZoTrFoW76vm55TCA325d4phpR2ePDGebmz
42Xcc/+612dpuudacTEzaimlVhFZCI66XIqFugl8uXnKBqn+0r4UWrqnRUMKr9nt
vE0CJL2mjxDppMyjRE1ac0w4W3jqgS3oVKhuLVJ2tkpmLHC0MvwdZF0SP7iLlQ33
0ZFHqlKIILQtwbHeNAi4cH/58jFwq3M1OXV5HjEJfzvdXbavuHuy+f4zOEnJKG1c
oK0yxxmFS1HXPcCGbm9mAyGZCwGpbBc4oTglgsLE3pOgjZbo4xDnvHfvdMU01Hrx
5HYCHQJOLvv+2xL5prXDJ2YiVlkrPnbwRXEJVYu4+BF+acN9jH/JYY9bICMHydXI
TK2pg6tqFHURDYPd+0txvcYGCNoWGQ4EucFXfcA/kyKUOwhSJfGDUSSfGLvAn0LB
ZrG0FGGy9O1CWbJMrqERDn9mueAXubr7SGgMVB1sP+lLi6h6RDuO4alaYECwIXGh
uZxfB8+LMug/66w5P+vJzkhHsxuj/RhXr+mm92fTWmP6vGjWr4xlsCrt6hq/oKZr
+fR+vLkkNwG6iaMi2wizAssstBo7QxZ1WB+uPy+tZ6SK/Icj/2zkLTtbf/FKOiFr
8jcvKvhYF93Zjiq/U+MPtpeymYV6JaCChXOLr1gexReYp2Q9C4FV3uldv474K8Uh
SyJlRdOKSWpj08dwLjV5FRe/kZ4XCvaAzPFs2TmQk9b0J2UO+cUOjjJ6AaHuuQd+
NYHj9Ku/SuxqKgMjjsWR9VhEw3G/bCUHmv98ElaOa6xDoLFChWW4ROdGmoAt6MkF
1H8KvpAVeQZwds6gCGBWlP/k9e7pg0qGqcI3euGjALHV8gka60Z0r/6gcOr0Nmja
+3Ttj1sTkCD7rVMdhiJgPZ4a66eb1uPRI2cQBiGqjoBdPY+8fHyVRUx/wImd/XZV
eGx468EPeIaPS1tSVtSBDtJ00b2OC0E4JkvSflYpRGCiTVg6j44BqTzqD2s5bVOm
kRTozHzy/vnC2lSkFN8+FTDzRs7Hpn6xNOMasKcCyq9daeIapxMIPujfDQsNkE1q
/pviwDx4vHozGBPEaiv+6OlyewQHJhZU3Dj6MtvzALqvxI/rd+ISsfPDKq4zLRU3
BpMHBAWcKpvCuUN8jfZCJJBYbJ+peVEa2dZm9mxawYDnhcZbc7ckugi+6HDZUL9i
4SF6CPxio8baYViKmdULZEzkLZzLjQus40ZGHJIve8fCNiDNwKvQKHl6NCmgD9V/
0LUncAaQ1WZ6ps0slZ+XZPORJaSr9CjXCpQ69nvQJ60O+9s/XkanTJZPNU1FbTvT
f9tr0y96gSMRNlM/SZu6krnANN7qGV+4WM+kgrKtWjH7Biib62pwzJkkfzvvR8VK
jc/SW2gS+77+xYQ/Tq2m5b+FgD8ADtk2EstYv5I+LsivFr0s0hhQ801Cj1PeXQfQ
crClCA/Kg2JrbqNvVEtQ3m0t8L9qkfeNimLTxpCk0cuu1P+pPy+ngDw6cyH0cBY1
pPRhGliA9i+zrfEvshOmpjo58J+J1isP6GEpECrviI/19dHnershbfFEMS7awmUm
n6c/eEIWEqoLD5yMiH/Q7wrPQpWolxRn3ZYiab8iKRElWG1hsjrDy/dLhqBclst6
bD22TXr5KKO2PiK5urnABratfoaFqMOcVUZ8hBRLbfH3CsgDSBkj0dFkDBlUFEri
bWre6dXMbQeI0eoKXvLEZfuAizMs+tWlR9IdrAuigH7xUua8K/yLyXKW9jMRjYjN
+es8OKcuW91/WsRF8uK8ZisI43HLi+BudM8Jf98q+jxJ19bDUwvVQ4Xvr+SlRgLv
yhE1Xj4SjeWIHDFP4rbe5CgfnnR+HAONlwQrzSlAO88YYMbNR7KoA9BSVuMoGv4I
2wriWtHT6r42PAJ/PeF37J9zKcDZaj2L0Kifxx+WWgGVThRHAiIlK5Acdxkmx4d2
vWih9/05wDpvZYWbVJ22GNhN/0jIUJZ/szqz66F2dOR1OlP2jhx7sMPxjaonSwgK
KT+XICkA20BocwvELYXIyd4+Xokf5LNgPzE1jeS1BykWfvPsF0r6rTp7ylg+Y+D1
sAlvnSrFi/oWDdsGPOAPUdFTyQtCqxRTpbMDMSInnhmUzz8GcHZeqNOu5r5Dmt/Z
+IdP1GL8UoQi8nq8GfYPSyjDDGESPoybcr+QZd+8uIcs3BZ0pX6Nu0cP1MAMGpQM
VXRI+W+05zLn2PxFCkBxc9TjJWUjFUJ+LaPLgKaykjxt2KY2gnKnXZoE5pv+vFrU
v51Hd6C8wzziWoFTJPDJbiTMWrnHOQkuYgCujUw0Zj2nblYlZQPYLC6cmvIiVYSY
6MSttA9Op9gAORH/KDVTVy14NtG+r/i4FKk1qsTqant9OJudhA/XzAEAqhslzC96
3Ivo70YfqOgnD3rkDrvKdDZE37CiEtu/ImttJEqtGXk228Mo7TdUpW1+he9XKZ/N
RBSwb2hS2RWqpv8W+RjSQIg5Cy9NfqFijEtJ/snYgwcirmkMBhF7nssNtlP8dgTk
f/Ms+98KvhId4G/ZpW+uPedPQkx/AFmJ/yO8PaOaPD4jG47YYmeMwOe2Gjhs+kbh
5NKTa+8hzNnbZAebBCAvSuVYHm6Ibiw6TarVS/UJJIAVIrcF8MlzlWKkE7AxC0E4
E5nbn8Cir2hMVhl0Up3aQE2PWJiPpY/rLCYdBkzHyGzHRdP5iRIT4p6TZuW9rRsn
6B0N8BaaAffrqvl7WomBAnPrCyaCkM1UeI17U/sLn7lTPXC7+ZO7FG566b0Yy4WU
4y7gXV0CG2BgxC1XiX/ETvYc1TM0k4qq2uEPgvfnBXoJbLeEe3la1Nx9z9chxOaX
w3uQZL7QBFE/PhBixuaJcJM6SzbxviqHlbrjJN0HMhuSoREoUHVquBZb+x7Nb6J8
TVas2ZPBm/eKguiBHG7Z8+NWtcFu36ghJmz4xirGqmgMNGM/aK+XEubUIiXaRbBL
sfrK35CLdItv6seFP/N9Svj7U7w6swphRec+hG5NQXPM7em12MwWGcNLBVXkMuLb
eIBI2qsVW55czMZ1aBd5A9b2NvU1Olw29BZzyO1W9GDV04UnaumIrdOMGL6d9+QV
x3au3FKBycuCi2D4FcMvAvCOMFbCiFuTeER7VM58sdbBjQHNIVNcbIe9bVLNHmiA
nM9CdRyx7NPQjM6ep3YbG4Ay2H0dCN1ueiTVdbvjj0mRvVEzA9IDz52F7QAEArNy
UzKxDopmSKny3IoOGVKugXdB11DYjeEGkiytCD48CGQfK+FHvXLNO3qBX7QhwkiJ
`pragma protect end_protected
