// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 01:23:51 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l0CG6jBmxmfy/6gkMSEao8KBT6Uw8zknx7ea6bMQfKWmw5ZDNLd2sKkvR14DsoAi
e1g6dSHaT4bDpmmhDC4cDvQyV3It3OYsV7LiOwkH7RQ8NgBXcJOaBfBvjjy+ur7h
GkL0RdOfMeljZ/GwbqXJwlQwiTl5AJyqVGLjI9Uceqw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5680)
wAFZn7J5wYraZ6/L/N1Jw1nwny8WUcO5WOmigm4kwun0pJVOzPrvS5IovfRskD3+
vi4BftXPMhPujAE11K4MGOTHzuMJVxD0vD3VZedVAcAJ7yYev1rxV2mrzLkcItO3
Icltg4rnlnVW7qoo8BbO0AELCyennOpCYqhzgqc/k4NOJ35lSQD8nBnAIAibDS9Z
lB5diyyf59nP2DRSmOdKmCzLr79mnQEZvZzvyqkSvdBpGQxAE1gx3FOQpJciKraz
HZ+tCI0D4MgCAeDzrwyx+G/+BHnaaRQAa8RGGGARr9SlovHzRJIMWEs44hCkInez
9zheco1ayjAAsc6IIV/d3xX57V8l4H6oNSh75QciEJfcHaWxbxKNj4er3DLSQQJu
UVz8NxnK0apINLtdBC8Z37U/hRsCQczjwd+pSJHfxQ3SwF0n/gyLXClhdkbLlczw
FQJKKk1BmZzdxOEBgZRMRE0/puDww0lQQiHY4sHbL1h6qiaz2BKLlzd+bVH3RjXB
4UmP2PdrKm/Z1+mexEdXUeruJnItAU5+HisBUeYyv6ivBqM74SX4b97CPikQLaqV
TaAfZM4t8gjlfTI4ZQnxvAtczYDzz/QAv3xxd0XnUUY2p6H2uIVSk0ARfG3Zp8O8
lC2KdGzKHXskcN0OZ1IL24BYQAWBxZuhagGTDZKkOD3eXpbvjn6YtSpEvsUvC1qz
3jYUkS1yFb83HdfUfjW+yi21EvONlz5/DCRG+fAL3UxOVv1vyAFSEJbK5v6n9eTn
mM6rLzz9IapgfK1yNNvAkmAQlQUlU1JqqSi6AZgrw8SzkQNAATaNWXpwl1KmThX8
5fR9/ZWBxWTtmpwCc3ROIhapPzddkx8hER9CK36g0/BpjiLDoSJ1hDRaB3lP8JsV
APDDX1O/7eTf3Qm6be9SbM58y2LnJwZUXSN5OroA9TWDv2YeDhbkH0OisErbamO/
zVmolrYvYPmeWaTCG8JEODl99q+hYHcAPzjJ2kz7rDKsserWR9iiX+ZVa2sEOrZN
zX6FBCwA9xoYwdaKiAl5L4WdWjc5frC2i+1FXweGHAZ+WGVwlY22Q8tzyJWen7Gu
DkxD/vjTjAAOc7MccbXKRsCAGfStb9/NEu4Kr30LiREJbAWhuHpgZxWkibt36zoo
FWQbpYRvmAdA4P7vXny0I7W7JhlI0VI67YqPXD2PRRfgvJCWsn7c40XD2uk1HEvg
5dDXkqO2eEwjH3xWVZO5PkNFKevG4oga7Fz20iT664lXNRc2tfAax+AsuJjJ+img
Dubjoi3eWID4po/Slf09gdHCIK24gJdXDWlK8fzTcGuYyoLDbU2g6qejcnKPa6w7
ClkxjOTFJ50ZZYZzlhLu5IZqe4G+sUiXDDgz9o8Qcf5mizua+DYbJxZynhsDyafN
1ygI7UqEpMQEdkOFQNukuVPJj82FxIvKvl/ETj6KO9Y5AHBlJlnf7PofeeYbn3ml
cUxCVIrMUlJzMbz9QmelHgzBIw0HE96pKqATQ+CIMl2wdizCimCkwPBeaLGKn3i2
BymLZQ7+UYnaDGLmTYzsIri5PmhfYg93qahE9mU5Dup4SMxNdQRNK3IX+EShd55g
f90dB4EvJDWSb3pCsDiv/DGyJWxahiR4EBrfyDszdu/BQFhtfWqcWu2fWjMDPKPS
1vfeMC0tTxJN4aub1KHB8WJ06PWauDqFgFgo1VXzUbY9gDTdJh+9pDd5svzuuI8M
IlAlVPAzE46taFI7Qq/giKHvkyAp4+C8sud3xH2Znm4wdnkS6fhWKs+mki7GaiL+
2M05Ztb5GplUHlZQF4JT8FGQum9P6+9YgfzbKTPJBxN3uRxr5HzHl1sspOO8suao
poThrGKGavMJ4kvi1yxJto8WvJ/Z2gCMBVpsqu/pku4LDDIuK2nGtnjjRW1wBqss
AAm8eOJQ+ltXDKJS48hzUdWiVrUiIyKT53jFIMuIaIRwhL4l7gEkMsUNvaOZ+1oD
vJ2/9dZE8e5NEL14UR841L5kMu3g5qnRHCgXOdvYRHqKHl7m1hI0D+rCAXN6RqYC
iwGzpKy0TbFLVbAlPOwubtc7nNUGP3rbd2xP+xCJsUC0Zw1DHV9Pa0zNuzUNhWIp
0dCYUY2YNSgIcJdJhDlgarMigmV4gR+88jtcBNq4atK1GBeQMiWLKKcHVjaHJw1B
2IXJUERvXgKMXym9gTPwohf/lHessrN6mITikq12al6oPBE8iwZG0UZ/9R13/l5m
sODY7faucmUwPIZfk7NTJMy64TmqELTmf2aY9NkrCU3wzynG8yQO1AwG/c1tABwM
L4parEVKqYV72DXXo5rOAHhsyRKassrASebRcNaKKouNixJ4FhTfRVvjR4K39zu7
NQuIujiSezjYoQDHDkSdrzVNsmf7G46n/B+1IqPnt9E+NrmQCVtcKuZVOZt6QroN
gFWHJhxWHvI+T5KpUkYEHL/LhLA0u2FwV3RpI8Q4/lHHFPR9s7wMZEdQqwHXwIjG
anbcFNNfH6dc09vdQIz+8jfuCBy54JyBG1K6lBR8oXcnJeZOK7ylT9uGnZF5tRTC
iphismVxN+qclHOrC65npFG+DhWGC64alPPsQwlnpuVh95htZPIrshPZm0jmLBRb
vjnFqNZIyXU/iqFxygArQhpZDJFfpk6TD6bWXlr/w88sICuaxCWTx+unvzXJ9pSp
a4e4jI+9MWdLIHB9KfnRJHSXAeYTYMNeCb6l8Vu2VAR8cK+U/sZ4QtJ4AlXHmosC
I6GDkPNQu5ABqCBbYJO9dU+e4bLWXpiVUD5wdpPT7hBr31tGKH+Rkg1iD2+GdSxJ
iVSXIoMARW80C3xR7IuhRn7R3REM3TAKQzqI3hZRMJIgzJvQoUv8XQhznPkL8Fum
9MfeqxbTc1dXf+f3HRJCvmiOUBAHIAsR9TNM6SEfwIKaSu05Bv1rNz7NGmzVAf1f
wm6CTPxAlCuA+ldSSKaZe4obkwTugnmFYYqbzgYYIAWOZ6XIkfHcMEFvfWsl5VST
9pBnCJyEH72oLWMk/dRB4pG7GMcGFL+Qkz4jY7DDFfR7ucl5IgMHXIb7MEdAeWs8
POtnTsp/rUzW3nBuYjC/wSROqhb5LNMY+AD8xGAeOaDDWJzKmxYj/MCs4PoLFCo9
U9zztD2upwDzPqR7Qa5ejd05MpYpxG75e3F80PFmGJK/Zza+NNLumM44acRNSST8
xa+XSPQSJza+hde9y8x65mp5MiO/AiPXbIfLJeemo+xmTVfV+vuSqzXuUFABLu8P
ifztFOdAnuk3/nXCJG1xbruqh1C7TdyF/yShAo8kKutNRA/hcSOXGeWuNKZRrmLI
HybEb3WiTnZpd/e+EzjJg3LIQ+xh4MzPdjRPbVXKB/gPXivHabk4H5/S7W9HYGj+
h+IfSNkq+aXXp82MI4z44UM4GacUIiTrc8mGErmgp2zxUiu1y5zfcKmVfHXwiACF
LQnIFjw0xBQjpSGv2y4kjrKocjf2boxZBTv3XIiNfoC8z49DpOt2+RZgmmlAbGnd
8EEp8z+8bpDKVliorq3CzXvwTdoFciHqt0pvBzwdj2tOeyX5kJYLKb99o6g6df4x
6H3+SuXRdFIgmGbB/8WVEC43LmhqWJOAILKJb+4NogEH9edA1x8l7e9f4yqbFHzD
XU5hx/XfOsXmTIPedlIzpW4b6AjCfZ9E5A+9hHCuRyF5KOlkSXKSWyNEsiuNhgNu
W0hTdiZhURAqeDryyPmnnrtXWuGDy7dgI/t8OrI93wNlpJoMJ88zCKxwRwRaASpK
SyD4IComiPXFxyaeo5aBWFGvg0FWJXXJsKV8TsUL1n4Ncoa9z0QNLjXvyHHKbVxm
CJbTABOeni4lvTv4foYipiDkYwNOSby1qkpgs4+SIjiVrsocTe0ULqlogoELxQ8W
71oSiAjBlTD6U9Hf8f0u8Cf0nOr2Xq+aR18iQgQ7veGWb+5QAkLKFbvs/MT5WBNs
y+m+Kz8Q83pMQllvrXXyTcYLbYGRDEJ4PF3CNLcKQez5g2KF7kcyX/4H/KRPfhn2
g6lpvCQ2BXPvIu7LOF/Vz2OZQWIxl58eDwOlwJzOunN+r9F6KMJQssAdnQ6z6S3u
ga8t6i167bn5AC9arXLg4nkvdLP1FCdGxFb3DDS/lVg0CLC5cTSpH3r6ooL029mR
WWDVUACNCUOcD0c4Y5pEKglyTIpRg28CymnhhsTUMxrUc9mwEu9A6WSbIQxW9kHr
vlav3ouDyj5L+N+sqBM/vEBDSE8R1MoqRZphIuNSYt6NJ3vML2wZ7qBqcsdXvI5k
cvWUeqGltJnts/Cnd+FYQ6CleJoeziz1WQFTJGN/UXYnn1Khw3DG1gwOzgfkCnPh
pDcf5saCPNiel4iETipmGiRRZwtvfbuszU7Aa/eG1HC8cn2rcXrVu9uyu47q4Uh1
QzApu+Pq9SnGxYyB+WT7zi+yja0tR1IWTOqxpnzdmDjs/7LD5NgiIzBoeTzHCbtb
OhqDZEJ4l33hJ+aaUocmQZyWOB2dm7OyMYgyiBBKVo3nG6KSk1og9bjYqyOsavvj
Nipy2kO2NDd+nfnPHGJmzldxxs/nX130FlQE1N91yg8FfUBSbpAzGAh15nwXqLzb
FI05hcuPJ6WYfONcAFH+CjPPu6ubmEEkg0CFybYVaoqlBxE39qAVWbIbYqfcpEsj
kWT9nWB+QpJuLgQhBoA7qi6a0sqXTiGNc+j+mgGLyIyWT68k4BUdRPVJ+eNIadP0
Lg35sBE974AElC/jSUkTt0IG+gIQnce2qpuA6Oc6MyBk077hTCK1gBbDO/yJYuTo
6Km2+0oHdAdshiRMP5AWXi9ctP8PNeiJnAfzfE3HcJoOMzT5kIF/6rdzVrfswwll
zuuuRCgVE+xoSJTkZsE3Km4M4E/vNAMcCNSoeGcA/0GuY7f/cZUZPaxVVprVl5CA
4STHowKvlsPNE55WyYmRuECaUHuvVAxNQYG58VQkpCiqxzlXNdVbOaygTqoJaDvM
jgAgtRcjN9JMmo4FUkFziLcrz58d7ts5X0cRaESQ51UtszyZ/8AIADK+Oe2iGMWB
HaWBShQYTuTbYM0M/q7H7D4L9u13OQ7YmP2gT1CdDG2FZSI9pbAnrk5uPeGMx3sm
YrNGWt0/uoqdZ1q3GXlb8zBnxzk/Ic0WFnaKi/haSDIYNfVeC79ncRO14YwdCuFF
OPByBh5NJ7X7K6Oty3HHllevFPQ5gfFGndMDUVZDQ+rZm6jfOg/QweVarq6ZJTwS
sNfagQjvdfyIq7HkSqTVEQzeRGtm1sS85hUn91F5DV2Qd6WhtbjhQ/cjlAzbPBnY
9iB+4//7ZjVBD9I6iGZCiS1yh+KIWgtlzpQVXYC8nFa0l055Gaa5ZVTE1yBdC51Y
HQerkifBSOXK34A/T3M8LByvzppK4f9J60t46JSPFx+lmGG/dgC8V+1CowkME04q
PeTZ466kpH9eO6eHX7nC9Gc7ulxVAVvAVoJ9L4nMLZrCXCO8hRq7JF6NHe+3cvzb
BHNQ0x8Mn9OyTwFg3ugR8BK7u2f6HHjv0XWw2HjTIFmpB202jMzEJc/TPARm+9+K
EvCO/4WKIhjFBeB6qkE8pvrBTz5SJSRpRl58OtHsJhq/yhyyKwAf4kz3XGQTPzRM
MJ4aN6MP/kK+7K6npz1gim2dokvEDm/qPVDreadG1SUsnqVMm5CgjI6oNVWnQu7S
Z/H780Zxx+bYR+VlaIFsmy2xEd30kbJ30gPOoA67DRXhJZIum53XG7SMfvfBzZpJ
g9qgQIJ1g9X4e/UHQOYsrxGX5XbdsTVg8N43ilCAZW3tOYmjXz9HjpHVL9XZ48Bb
24h00rBFd4gqj1CoxPAOYQhxOuhRSVrv7Sed/SKDuHeuU2meOeRL2SQStWqSDfkM
56OAdEkKrIkh+XX5XyUkbovSLWpUaSiqHVMXsaUVqeMmOlTMmY4uaGWeS4DC3dUU
HWejasWo35vl07o9OYjgsBnfF+9xxOxMN6SMATOZwkvnLDO9cIiYNOfPBrVO1pGO
LlbSOmu6To1Wk7QvTvqL5rhsVUtvbNDGtW5i7fHGdSmcD30BzxsiZ+z01mgSC3AI
JyP6LoVzR9JUnjxZ+CTbJG2YFi8NnR2f1QYcB81Qomt7XppNcb6joofRfrXWXNBi
pAuNCQIECbFI5KK6LozTzBvwFxseYVwRu2E0MX3fu6yVoBvtsFK8UwiBqkdoQcU0
knKqOrpnHrEsA/nuVoy0lc/gZ57blMjp8PYT9isx8qh6oaBbiualaVXORktrXQob
eZQr2I9DTK9kLsK9bgGow59ITBK3onWEYac0k35UxWNxQI0bxh5Fy/O4pYw3yPJE
q07MmNFb3p4UmBNCI2MQDS0b4vGwvQDT7NRY7ZOBeVyJHOg6p8FGybRJE3LFzkFQ
QaHe3ZTQzlVe7nm7jUjQENdu+y4yNxdZmc1NpqGC7TGU5oN9xkHdOQ5wZiioKVnu
YSASu04OnZuItkHPf4gU47KnLk86awbO99pylnXP7WB4gqjMULc/oIHb1otHwQcd
AkZhbUkdgcY/4gVw6mF7TXPt2Tb5GyP8YRfmPlSSy52nGURq7uumT0wytX/CPccx
DuJhn5AgCaH5/1clq/C1uJIzVuujAha+qr3zDZ/IfZONTPdS3F5sGEOyjTojUZf7
LuFuHeEISlui2rTIQAtbjlJKp+5b34u1pmwWKFL2O8Wn3OatloVybNMEwgyEtbd4
gLjOkNXJWzsKxpMst1F5k6GiLXMxRUW1HfVPgybWJ0UwmpM4OkfM8zciW8MMyzuQ
yhRyqr0kMl6Gsfic4yfrkZJZ33a2aVPYcqdRPTSKKHeNmstsvszMacj1j3Lruc2v
da8m1P+ZlsZcj4bo6ChhCe0FhexJfobo+NYv1135jcjcQ6Ky/N9oOV2YaOdwpwle
AQG94s/huTXxawsfJg9t1eiYqtu1je5E7rJcVOaivV2w4Ol0SDh/rwHEtjxrmzdg
0a9Fw+urHoqICTuB85SfcltV4VfN7hclUbT9Q6rtOJrjFMa8xR6+b1WpzC1dg6bE
tYrV3/mXfFlMcEygEadA8NvWdRdxlNnpWR4QXsqLpun4gCHaA7SNl+6t78GRDUKv
huF54o63r3NN4+DQ8XPx8uDa7btnXbetaGqJNvlvDpALQfenR8MPTCeMKEiGoU7f
PYBSCKq/Xt6dFpf7N/aALQqMB0yfYXi3wvBPhhxc/exbE+nVjEo3Z3i+XHyzslSx
c8FaGIWcU2WEekRZ8EVoAi6yqMCHROia1jOAbjzVfN72xjOyvB5WBMgTc/+JqIeU
XKSyh4U9hPH3tU1hiM/4VFpy8JPyO9EnK3tCF3v9HimuSLurNwFS2OhWutSWsnZh
s6wSjnUee13ZaZXagDeBYAs3spaWiYXAXCr6bDmFt8WeT/shxLx5i9QBNZJ3hYL/
OeqERIizkN4qyvd1fn01yrjuo1RCQmzYQFcJhMyDQy0KDhiQ01BTazXmLllVYWPy
qewlwR3tp/ue7OCthEWDQ1RvPS32UbHleH8hZbNwr7rxbtc03tcjj4wplI6t33LD
Uw21nSe0HKn7Afk2sIFe6w==
`pragma protect end_protected
