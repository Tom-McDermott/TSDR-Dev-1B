//__ACDS_USER_COMMENT__ (C) 2001-2020 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
//__ACDS_USER_COMMENT__ ACDS 20.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
5m4YHUczf5Cjg7T0Sd7aG678cSHbqV5SSoZzwCYse4CX9ZDRF7f7q/OQqZ8Hsm7v
1qe5P7ikTaZzEdRXbxXRV8XRn3maGkbanTZXREbrvtkr2Oa9s1P6YV3MJ3iG2yrd
rGGJk97ajZGob0LPpZcaJfioQJNNkHJ71mZh+ifo2qkKWg9u+192rg==
//pragma protect end_key_block
//pragma protect digest_block
v+v0o8tDZXE8AbZNyJaPab8HN8Q=
//pragma protect end_digest_block
//pragma protect data_block
lTWhrZSKSTxhEVeGz7a2aXZT7tYvCmzy10IvSflSO6xcCaCXFHEKO+DuctI7RH4m
pY6RBX2e7MqmtCUP6YwDXEn8OMAGQRZebaumCKYbIgbzbVGB/SARcikyEBtRyksA
0N+3iQfwVVWB0cY4TEJExT2muhsdY5hf0E5P/HSoBrjGNWwdX6Uvd41TXgGkBevn
1EeRP4bctkGWDhFfAI9psJ0MWijg2c5Kg4XF8inFyJo19uEn7gbCfybbmgBDDkhI
p4hfQ/GhPtc5nVl6XXdX/j1XV5FHBF6Pw0rpPGd1nwha6DBQJpyzAjvhWAsqzHLc
oyHK9oG4lZJvlDQVyJF1TGj/iPNhkhSlcmnj6/5yW/QjSyEwbU8HtFc/sxAaLejQ
Tz5rKu1u3EMYLuy7urCnXAEvnEKEpt20dhKrgYCPkphaO1Dnx7ka6UQGeniDrBzC
fYSEWKzKj4ZgQBUQGjTUJ1jYsq21RTjdi38UZKwnOBfbL8VQqKd/O18NiL2MFoXw
YlweTgkx2OPlRXtPEInVQGyILE7LqPd5SEHgB1cRkteZpZlukJPNo0ZYTN11I+PJ
/nNCkejeBBBZ+uLQaK2PiRUQMDjNBXF+R/Sbb+MDFnAfL02udzDazPmZkauKECq/
iIJGEPmgww/hOlTP/TOs1qj0MoZwuH4B3LpS4CvwZJIU4b8XmMPYyAH2m39TzkML
dyDebYMVMuc5QwBNH1SWvq+KBOQ9NSVTbD8b6MbX1INerRgr4wFyVXJwajVWHL1y
wEaumXfynEKAQiPLSst9fcgmp4lwKO1LhKEwgHM8CjIpILIHo3CCuWMKuS0oroUL
GFfHqKcFtKbsEVtxWWSSWNuRfhbon7qoVowLC2cgdNBIikk9MngMjaKNGWHDowTt
+/EM9XCdOZ8AwVjO2HWNYmJ71Ec/IaJYnxAr+DCdHOKseW+B/galTBq2cTLbGZHU
96yHWP4mCHhfa5AAdhN3ElCPy1fMzELz1XjulKLiTooR53nbZPqdxcVkN5yeGFxS
jEdhX/dSwVVYfwK/84m2isnOAkaH6w57b9bIklc2D1Z5msxwD4CpGhSifkk7TcfH
LM+4djYu928JMzg8CevJa5LlxVbu6YTWAThKP4q2JOxeEyldKVcuynbIbc6Ttbt9
Cdz2WJizOD/cuU++kCW6WGcau+65GTSkTrdPzK6cghpK1waZZ2Xwi6TKeT8I5JDA
huotWJ3sVhezcYLrDnBKy3z9CAhGuwxGf8IOoXJBFMbY6TXFPnhmVzoexet2hAdF
3pCSAECdLL7Ygcm+2R5k2w6jXKvskUOhszWGM8mI3dQhfAxeOSO0XwHCUNKwU7UB
1zVaQCNYjdkNpUpAbOczUxmy67K5e6EabOrhpFZLtxT93DZ8cusD7dxQP+wNtmJk
1LuTUj1obUcJw4K30Cdx/+8I8bx9E53wOIjmZWoFxuOGChQ6CjanjUhUUQAfZP0U
1ipCo6lw+6paDfSTUgBScSl1qsNfP1NxDo2ezvZnpGbhRPWWBabiv6o6MHbTMy6c
1OYPdc9C2z57mt/92umvzIKWgrYo69LHk99AVlpWL+uJOCz3FcN84IHnQpdkYHQW
4aaU+lFRYyH9eES8qR8NHmDqSTslu8AMJ4D3Ax+ZF95pUgsRFGZhJfgCv5/pUTis
n/VJL71r8+eVyiB5loHljie3lnLPrKn0+Ik2oElmV7MTVf502oFSWR4JTKVCc97t
f6k73XJGxNNWEHYwPxuGsJDzuDPNMYez4Ls9rxfvilv/oJs+soTaYNXNefxbMIgD
SUKsP7ZzuiwMWn5+SPTtWHaWJAt3I4fJde6L7OytKX1GGoKnlaKzJKL8BkQQBSZK
hsS9PdNHSfW+rlaW/LuGPVmMonGon04C1lOTBwbAdrOWnWlqZejx8nQm641Xjzis
ub0xrQf0XzBN2E9cBcHrDiZQqEVkhO0ng4RNrYvnvczKEduBbNAYenVOknz371L2
TxsIhFvEQ1VG14oR2aENzJ8NlMrlP9paMtlSXv/Zhmslcb4AMGfKTjAc0rFRyqzF
pjwHRzDxs0Cf7IvgYgoz9ZrqY/r7E3/JG4XWF3aiR3oBbAZ0W+Aiwz7mhHCuq9Db
V4KiTwzIquBPqpaUQHS6ND0enn4ModxTZMvFmsWuEzhAph4v2NSMPUV/+592HnVh
CFwvv/p88D+/HVcmKSQxnq67P4vfWMdmRAi/qWk4Wf7d5lA0qRYTYZX/XwHBXW8W
2eUksxg+cl6HThI0CslM0+YeQYPwzmNNhMgh5Unn6RKS/w0vpb6BidcXZd7qtN0W
HTul3o25bDWRzubIzGlae+824CPispRNlJuNFI7uPiy00tSMN8WUV+P7OoMLuL50
7Xh6NaTyPEsWfg5IywPbMAONexwdsApop4HZZFjf56/vwvXYIZ2XAddzoaCfozPI
o97meufnz4ufX4YM+3gNpslLwos3afmsZKVz2VVNt5ngP26Wsl2AfyBzX5ZV0T+K
tlMmIIkpscMpDvb0RMHgXTY/PDw/eND5/PMBaXpNnhvEr9lmfVS14En35eWWsaq6
4yj3k9CJ4eEPYFp5w4cssFIMr8K4B/ie5g1+jKzyi4L9Mq3QUThEKBVkQ3Gs4cI8
i7uizN/12r4ghQtPBz+xxa8aGZPcfTmB1dHrdQ3sid/DY/aMMmZQ+MiV3J7HPqTd
nLZlKLal7RCfYg8odNzyurar3gxbWlC1i+0PibU4qdVcMwwZmW0DrDR3Pu7ETCW2
SkOcCgvG2e6mbdxcRkZmBmzWm+129fTyIfjlWslmGn3eCC0LTUWrgaf6bO2CPfxD
EndkjuA0ZmR9JOKFrDUo6z8zRwb5xsYb5PAWkcbh1LFVgtTO6+CXEYyW9XQ+XVDa
filhu2qdfIV6mVcAISOSQckmO5foGKmWHsPFNhNL3WxjkgJILdyLO+gb1Cu3e6kn
7y8hddoysqpHfjaMG4jRaZ6G07/ZGBzMgHjsqQXegUWwhVfOz6OdEVqprxdbOkmB
q1Hg5/+bbEMCt0HweYldTUKj1ju+PWy+aXOiSMYlFjUDTCmF4M1oUer6g/u15Qqu
h8cEfgTyFJNI4mx7zm0VRDGwte/+QvDaI9EfzmAuxUM38/ixqv4blYkOPgISeAmp
ZoyP8gKcgYhiYX+FLpPpvceRfdiD1xjIZ5r8ZYLeRwieJbsR9yniPUwo5UVezpwj
bbN4QOdFAMgnT4PbyV8BKWpAiQoT3jMSE20pkNVxXg6Fqw+fWsOYV3c/eqt+d2Vc
bY8FtJc9YFsI/q3ep8RXhIHHEo6tlhDshURsUSf5XSv2p0mLYkRQIIf92vJ+7h67
ZNTdr+zob0XliQVUdi45DX/ah9C4zk+kX3DHcKuZ/9tm3fXyekE85Q8hZCjfCPfr
Fj3N7eNfEB1q/0Nqrul+GWpuWYpbeR/ruWwzhl4LtetTlF8lglwpb2RwszuolWPP
6fThGYzMrtCH/hFtRYucGeU+Yzz8AkjV1QCD/ylssyXPSA5qSOUe3KxRs3zJXntl
ht9ybFzXhhf89TyhZ235BBIg2whAckzlza1cqMJynyWif8BP7vbpf8yJqzNkyiO8
pAcYMiA6/l+doedw97VIivVF7iODUV7hrdtkrGUuFy/iinLQlDOCJsaVq/zCvHz3
3gbtmoIakhTkozafkCjpiKI2vX4o5n+dlYaH+Mg8uP3E2+bMCCF8QEzRksynkl2X
jJdFbaWskFnJCCX1G8OYgBsIDb7NM9TvDicjEg7o0gRX/Z0nHF1EBMn7wawEN1Q1
2s0ZdlufuWrqYlGvk/w2k2njcpMczU7VsNCjKaNy4ervDuHvT0n5KAfDgsxbRjmI
mtPQ+Tl1p7OqSneV8sd+yjNu6fajN13Qqp99kG8C9Ynkc53Ofz8gBTqHAvAIC88t
M41pFRti93KON8+SHFMcgLrcZ7jNcvf7oIegRQy0QfBRvnVQkK5XK/ZAsE/NKIu5
wKqJz4NQ+Xpffj92qFbsBHpT3NQKM/426PST8YL9KH+CMJWaKKLjXdsdXYaFgW5C
hFypmJ83pIGGHsIzyxXc1sQVkSYGyVK0JeqHnQmVR/nx5VKvdEh0WR4UHIrqz5JI
1wdg6qV3tO/Q8trv2uj73y1BomxxAHYV1WuoYqbkucEHPfJ/kghnTrhhNDpX2njc
dH6qIad4FJ3+AMofDKsjMjvS5L2E99kFGE00/pDCMARxa2YLWy6gU+uMj2f1NB0k
IO93ijoj+m8D/poKu1HuW7YkuybOq+mPDmvr2X3U6yIi1X73vG3B4YUXZuVd+7nx
kXNkBCt8Q1EqYGy+i/iX1nPPhhW4VkX4pZy+CqTiy97MvgAQX0O/wPZEHVI1Ml3p
s+ZN1CK92D81XNzJv7gWdD8qIa6p5ZJcMwIY91UDFYxnq5VbTDLJn8ed/J+B/KSr
YsdDKQrCus+f+/uzba2EMhJTy6sjK7+XKUAxSjHvytPjBx/dY0EWAQ16FdsGC6tj
NH6bdIbAeWs117rfSsXI5kdSrZT7frXOvevmIeM2ZzR7J2OFOs3CPwsIE/7z83tc
GB8avJEf3NBC/hv7580oPPKSknOdA1fthINMcLziO+sN2FxpOBSpWI2YqbgKGr3/
XdNbZXkvSuHR3SlJXQafwkVdLB1CXGdDhs7O8wqATGMSkrIW7g2pIoukrpv62Oeb
wKUiTbFCfuvhi8muxWqFrLA691Rq6+alaFGEJJsKhkorVc2bTO9uVJvVH5u4u4ZU
ntynpKGO+K9DRVVMFuv75APKeqA7ajhRw3fcJZxvVPBNioTWE/O0vGa2EGcXgehT
UiBZ30rb6H+s+4yKI6NxJDLn75IkvP69ysI/q2CbI0JK/Tk0keEXVvsCJPQADg83
5aicNfsrB+YxAh3di440cqMQ5+Rjm7+37xFDs0U9Kpiv6GXn1vabpcBHJmMG5IdP
oLeKNSa7h0HGlgnvD3+15Q5b0G8h1lfAri/SRrphrxW/TvuiLjl8Jlr8lQHxv3bj
+pWyy5geJElMwTPI+Uje55Qp9oUwAMwYNdS/on70pM872j8s+pkPLLU5cYPUel8/
RP5wv/kGIrOJG4HLf1mUCWCJgSDms2Q6cGsekwh9wXyuPbWj+dihXPEJuuTQW+Lv
YniTEBb6Z9uw9hYWX1BTqO9EDy4sM6WmiMk5v2VeLq1x08CQTjqihqVqA+Nkb/d2
j6DIBisthMdjsylwS7oGHz/oJf3tcWM4OC+0sHRnxVqyopc6Zmw7v1hqeATklFle
PwNXZckPUj6LIde6BfXuLYnMAJdTsj9wXaRqhv4jtM7MhEsokooQ824Rn0/VJVb/
bIrGax6Kru6rkdI34ac6cvfv8GNyo3vetSiKcWu8SDVEfZ7LsWhQgEiOC7Crar/R
82xluEYwBCtS/8OK8U3HVDCrfMa+qBi73DSkh9fAI7X9a8TY7YhaE01IefReKigF
ocrQeFbUOJb2OX2F6wGYAOkDQ0u87NikohcuDDal54LXv4dXyns5LaJfyIBEQQaB
ar6VcySunS2/74IvqOTpCSsiPvL9XhrhotOHWClx4mjz9TfqSVXQ2D8xUxKagr8/
aqMUniE88OwOYQS/CDluxJflB3u3BNko7mYSp6tc/eqmbT6x9x8b6EcLT8NLKoOH
vcdKgOmZQoXIw7fYMiY9yKoZP5JPbLYAQqxgg0t7jyxoE92z8BmjsBhKWnkiF2qC
6c7YPcq+yBDxEIhZ7Bunv2uMdghCbUlAeF1QiUwrZ5Adk9uoS0bHanoVR29SMGVu
Wn1O5wQovw+A3+C52d//v1ytjxPyn/ctsHLIFVuGQnl7FUyetrHEVRz/i4F0mm9Y
Bl3NF1hlAU9NmhUOLzltrJEKw/mRWqaoQyi7UD+dsk1HyzCees360MCekA6P3eAN
9fZ8G4Ld2ZEX6fwca68iN444h3hes5JpQlXwgSHSEwAGmmlv88FvmVODzdphNgbR
Gb03OmZkfPWEmfNQNuDZiMQC24x9QjyMYPI6sE17JTu7nwoRNHv43y51zfMrJJaY
EClko96gh1+ijzv0OjcgF85KN7kyBEuppJoODbeKOI8MwbskIge7tcSf5c5k2iSS
iqwy39oIy1WnIuo1QDEJ0uj1Lq9uZnwLsCtq/AHZ4zfVuUqs+rhK9Co3cXaF5sL3
ZTt2sl7s8xFWjdtj7MllDMukuOqoQ0iul6K2gdya/onPH1g5GGXqnbLcl50Drpdo
BkxLfrX5A5bPBcCyZw+H+ZMMdRtaImeK0sxuwmmZDgndZYzZvf/Il73txHj2Hy1H
zm5vKOn0Q/4tFNPGG8HjXhO61V8x/OdXGeqdD+KPdo8ScMA0gPrhXVpLFbX3ZXG9
CHKdM7JXmo1NU1+VRiauYI5ayFj69dHE2na6kHosL7RDI1h1EGE3ru0LwsCYwXBt
xCubpgdhUNHRI/N+jThAGrhLwvjmHQUhU62Pwg+3oiygVwg+fhDtfQC/xLw5HfqR
9xIaE1Kedx8M/kjOhM3Jg5NC67fRlbWwmA28IkaFPxwhDaKPWkIGMwLf6MKbEdqU
wN4PqxlTRC9P4c22n5VxdY4Fk9/ZyiHyj7KX2NWd8FD6JdVTEKc0vnq+z1nDBLzE
1L+MOatjThwNsonlw0XwXCcaf71MJmXlpiKlBklAml1xthCc0cwij2E4eZC06QLX
UOLxz8c4y59uXVHXmBk+mFjklpcTtF+KxIBvvzMPS0d1SNgIiktCe03D72wymHrh
1HCltpHVnX7vqbMt6FrcbESq1XVRUbkahtV3H/qa3gWf/vW+FGLXcFy2Qf2ZszoC
ZPrdZtFXh8LSwsS5cCgg+nRV5hbJp6N3b92vg4YXV+/RCtDxqO/lSLnDXVp0AqDE
yy9EJEEJVye3CUvrlhq95AmdxNUSt7SF7omwp4S/zmYeUJFoqDraXA0nKGMys9I4
TEAFRdzHqHe7gwEpoeUKwrVra9+djlpErKQF3Z40Iog77daMIbeCb4RjDK3K1UZJ
2fh8dMDgOaIwo8XONvU+l8Ft1o4+esFo89TRLNJ2MxVo8BJMSL4bX4bkMxgETvSN
en0n6RpCc/+8cplAHc9HtcpMPtPnL0wAv6Omuoye+dCpn6uV4a7RLlGkCMCZtGid
Dt0NgsWU8Tdqqaz6YuTq4IUraeaP7SRQzTqvdKXyIrLNoJX7VMhWheeZIftvfoWF
l84mJpPJAQWIqbwnoW3ctY6EriSO9htZ+zBfyVimhaFdLWanmHw/SSSaHoV5sPd8
vbIcNbY0s4T3F+fHw40GkQKqD8W8aNuvP2PXvKbRVaOi5SU93BaGKNZenA7Breu4
o4qRDEY2BAilbryMs0lqRi7Hdanha2Uibe4unTps41LDL2LSwB+JlWC0zGjxuApP
VRP3PU9h8CfMKuccXMZHvOLnI33Sg410SO3v/j9NJpXLA6ybISyRVZYVw7U2O+nn
fvT3OELusQPTpCP7cFOQIw2/VTYHPQt9fLLP+7nCFrHsqeu6MNMlKeRO91egw+qY
ImQIwFDdbUaQoGHIQoqT+PfNHLbiPrwJ7odIm6PO2pumPSzCJ730BLb8nZKCM34D
YOPSoJRBfw2NjEX7O2D+eCSCiM8OPMjV7tlX2rLFF0IJdDzNOSZ1SkxAhSNuNAM4
noEZgRAaWNaXVxAwDiYFmix3oBm7AVWN7V88P/WdN+gI7Uc9CNlWhWZXWqTZCDRa
5YihpAKe3UsPPga4hYSPpWsCx+j6mIFYmab8R/3ijFXvPa3qXO0ZiZDd+d4YfqLa
UGW7EPbXBea+tlINa1iyQwD6///0xdSxRoVTG79SkTiBNiceVbf0raAqmQTZ1MQ6
ZVni9KbsQNX2LufAGmscYzHcGAsI9IUuDC2T28VNK6s+VPZ2szXFn4c69mW+OAei
QuNy8wgtkFD0Eb/ZsqMm+RI31urFgH6QaA6S8ZnSy2o1x6vcNcbFQfHQwabrILaZ
SYWg5j1smbka45iT6b/NGfijRdUTobDIRyomQPnfoHhy0/wU34tnNEif+kOMph+m
SekzEmM7RlpAt9YhWuE8plMpRNYvpru1WQaiEu2HQp3l2zR3WbAcROMMiywufDG7
Vo16T8i5QVeTN7nAHDpdlVUGJx98mBTa3ONTFGaiLQaGq53WkBSWNcw7YlKnzlDv
S7Wo+7bCCM76Lb+mLLals8lwojg7g8qMSwjF2B4IJHCkhRiJ7YA1PYo/lezNB+Fn
IulNHWB7BhhzWl/2aeGNJFQWLQqvjFFxIF1/TeXFflhoUsKhQBWouN02edSTUX79
dlCSxXpblrdCVshrKr1mEIKsrCgmpWYQTzJfbExdst8m2b78d5ZEEGF9wUlc/jJC
CC6xJdnTs9oFD6XNT3PCUMfT6NwdXT4UyYRMG1gH7eh6xgNJbxTRsA6VKaQ2Q8wr
ktXzbJiGaORnlqidKFZU6zGXhc4kWIYcsnUTp4jgaC2qTwhbF56lnT83s+6QdLP5
SjuiT2lBnobnM5Oo2GoCzjfBulIbqA7YwMr9wJYA1XKsbGP6W2mmtEMs/yT3zC4y
mWjCMrrXoZ34Ju0ELKsJkX0lcn9XjZxIOybvHyX9arnYaAm3HLdJs17NOcioZqTa
6xk+mdPGZXwIna2mcGbeMR6Lwe648iJ8mxp9PBk1Up0FOH4dzFPL8D8LrzZNxXrg
ePhVD4mqdEgSmUnefunYX0Bs0Yvq8fJK+eLMO8X+QdcNvUAt752HfT71AiF7gdI2
B07FDbpC45tgTInr+g4HRwXQB5fROxj54J6A14hqOj2RQVLvVS3FZ/NHSpAWUsT3
opbgHRdxfeiWVgWaqUWyISaQ8bE8Ik3Izs9dtMB9RKdlJZYuopInvxT3k7nIhs7C
lT+oNjef/S1lQ6LVW/JgyTMucBHEYmG2e3Me8/1mEgZMe6n56XaB/Ah4l4G4EMKI
klR1uFYRh+wJ6HFLL47aD+UUoY/E1eNzo4DsuZtfr0ZGpCwRw7dpEFoFWZk64yc/
IrjnrtNCwGgNIEGX2qmCkQqcEkZLbgqnXNjn84919bNCohxnmPVBORlkj6yA4kZY
+dDLGVR3A/Ex6INVdyL8VbvhdocZhH4xIQaKe+u8x89k4++QAQTHa0Kb7tOW7FAS
w4dY9xPPePCo/yUpn55gt7J2QeCVolU/iSlj94/8BGbErIw7/+xCBCFj+SJgd5aG
FkWHQ7QMCgiXWeaKnyrP+PASTLtgEhUJdbIMeWGAbVldyUF2ul11GQH4+ZYHj76q
GThgqaJ0GYJJ0IOc0nogZaGsSYpFF1igSF9GxphiMPD99yvi3FsQt2wBoLkyhSs1
dM4IXWj0QYOTnSDm0FswDZwMFHWA0RkH9qtBwApmEjY72gW89ar4E7UVKQqEAfE5
GbcKaocvvYuehPhnP9QlXM0h7AyjQ5ZmHVTjWmetKFpoKypZmLn7JzRWbl8ZJ2gY
WKZWpZH8sxMVib5fv3rqxdfNZI2VDqLPYl8aJvTuJfZT4P3xkinrz3w0w/L/wpCY
2DsxDNdZoieRy4s5AYBAtUcYnAqF8kYVQuq5fPJEaf29PrfJaDkBCcTXyCuWj/cY
vMDtO6tRNzbjtAfDKcXKufRNwHypyieS8tCbgWbFrMNRyM3IwupBOReLj72JVvrq
2kHTxvwZhD8x9eTLd/T9xinPcC8aj5h8YQY/DV2srYfYdg2vwWIPEyZLKh5F3m2I
UhBkZST22OXDie0abimSWcKFM6fz7BAVd3FZCkIJjCX79b0thR3XE5fO3jZt2LYv
xyZySAvafh+K7Q1AnURpYAZpi7wLKGbPuzqy2KAf37ncbMskYF7NKcenvikWQxZo
XmxIyHO+aTj2ZJ7lx6H/0REqGelidTLpSvafgobRdPZZ2nLlKGl352jstUGMcAP9
9f/mwOhyd90OQTgslvVu3ofcbQLD/B/cBCdKsXKpUH1MOLCBKL3An+v7A2uiyVAm
i4dza4dumZCMlD3IedBLi0PHUR2SKtDgWsKLwPqpX2IyYD6wwPz9znNT4FioqYI9
0bQnCJoIYvHNLMDiXymk16cYmOgW+3dRQXfZtPmVxpqTXowxFC7/6KFWS+l5ptc2
DpvVMhLHeqpb2AnMaXZvSOoMa/aiKIH0hQdISdfAIDK8Etp6pESrfWuxmy7S20mt
3NIoC4oRQQeu7NHLP98GWEYDWIy68wSJmX2+5lqZJvUnUsI7Z4yJBFJguCH5umxf
NOkknPTRFShC6R1XHQmhVa/+EA5GNrlbFN6oM8Hu5KEfdGgmOUPx7xYGbFRuvMug
TLL+u70dnHSt50Pn4ifG88NKMRryz4TllymqY5OYCnN6fqJ8z33m6jUme4B/xbe9
3BnbLN/oWOKHmFHU/YMtcRcHhe/x2bf0UtJor2W+sKvTi2XKwGBM+2to72njlfGI
MTYgOOrTsccU887blFjONFcaKLS05hBXRC04onLcUhxtr14/2Q1JoZpmpihTflA2
8IGdndfOYzB4i2Bmp7ppF/1a0R0p/FHiHGn/qZwXN5OUHdMoydYvVfeNFjQ6mKAu
fv7QIrGY5XNIJjoi0W3gCLqfmcjvV4NP+uoAQWq1NzbBJU5eqJIkRGckwz91ndX1
CcxfuTPrwmkkxlLRhAkbxrympZIx+dRD0Rdud0s0KnJrByBgHWlgaYyALnkqS5Bo
gLP84ccBpZX92bSu3XdFe3vQswomChsjOmHL2zbu4wD6PvkheOUfSr1xcTEJmhhs
y9BwNV2K/fEu/E0Q38Zpv8hkzompOkvluphdoM5Fi51Ipq7Vkq7FtP/HFQmXPGge
hE5UX7yxWYZhCLy2nB049ZkzPbXe4ofGMSBso2ZDD0Fbq4O4N5KsS8cnA/8rm2Pq
8bjVI+CZMcfhdopL1WWgJCqErGPhovmlLRyXG0kXNKOM+hQxolGGg6gH2UayeMEU
s7bbf5G0gC6EbiAvhKHzptssOrMJVscjksuSqvtNrlyWhScPzmJCf4iLnmJ5yV+9
cC0bZn7GntMwRf5mNQtSlRErnZoinIZVorq1rJ46tmLr4fio+2tDGsy78YJRm0i5
xUuO7y9BVOX54fvVtb3CjHpVjzFIQRdlCk5qXAsoN1VlfG0ME5JFjfuWk60itSaf
Q2ZDPbjPWUxOMKA954MUurrQp3ccTw+iNG7aaSuaTixxkCAedPMhJATfCDSzQf4Y
SH+zbNIiIuNoc/v/hZOjtLppaJB3ISktsw/A25288SdaYiwRSLolkER2qdsA2D9b
JagWAPUPP5D6AZvEAibNg81TDWtUJTLdmEOVXj9l6JI5or/nC62KbsKqMC1Ydlyn
0IFAZx5Z3G/IbDxJ7D+RG8rp0cJsuan0O67sZPWXptyVLiOOWGQhfYEIG4flCtnd
ERXj+hjw+yAYWDK08uZ0DTRU+D+VGMsIPZtXK3+zXT18wHu7xx9NLEOD6+gMw2Lt
9DbRlA4JkFrjqtv8zPuY1mu1n/z8Nn7eSvkblX7RPURSRKCKn7KlkPhqq5LS9btY
VdKlEiop8waA7D1i3BmhFhcLoUmGEImDJ7mFspn9kSmP5nRdxbZ5XH8TBivhi7n1
+TSLUGVJzU65tN3aMu0fAzEV+heXd5gVnWk8G/ygvc7qQmXU5ie25LffutLeGs1e
Md+0uFR+wWhhjhJSY6aRxtkTYWeQXxRcxO0F5aeKjvbd0w2aOythh3jb27s/PLxs
EOp9N4lQPTwrfOyhY3hI0tl3ijUt1i4kEFXfUTW26Dl9OmehfjkXg3k07mg74/xz
yyQpE+AfYk+h/WcLVB8Ud6kmYoVaWAX6El+dPPBlYwwSdSGAXX89teJMJFIU79Bi
JhUfn15vLsIAfGAKIi9J4PhPv4PVcnx1aLqUkpW+kYAv+iYouw4gWnC2kk7PC0Rm
mXD3UT9L6u8398TGtHT7otovDn77lCrxRkmgPEUagFxgbe9QTdhe56C4iEQLXBtS
axROATeLa+V1pvQ8lE8UpoJZo0KbA+712LGBo9qZNYMD3DLVcuUtr06UbOYPV2g0
HPTtLBUHI7Wn8dicTooT6tjZOiFj7vfcoTVNq4qDhRBQilSSJU0znBS+tCO7zj9Z
bURt95QzdUExpSpsOisEQ4sswGDpG0wpYUbNyUYRlqiarrr+wYb6zOck0O9sfnXq
1EU/zeMH0PA8IwEFYHjWOjXoZL5nRltYE0Vyo2zEA2Bl/rGKlnnSGtXCnNS3nHoo
88uRKL8HwfgD4LcZpfXpcwUtaeGbzmMBIUxO8FfPB2eQjR4RnKEAxqZWk3XpXfBs
bajU1Pomu2BlQVA8VnNPvDOj0lYh9FEcSyevxEVP87bKIECeAS4tOXsFz79nPqlo
NHFBz2YlEYaJfGQTys4bNRhjUYems67OoLBMSC7HSjfDhMXiGnkzGcQtWvLTeeVw
GWtke3IYCSWIBCzxVsWFbYmk7nY/RlbB7SFRKAWVFOVm3Mr6ae0xeLjVuG5778v7
rD0AD53rRwFa/i9kFGaVl1RRm/iiEnADUh00xKJgF81dNGfFbjlz9910gmwQFwdp
dlH95SKtECO/PWxJvfN2hOEtTm8v+7l7ZSg09pNMXEWN/XRLVPQMMTiZCHuAQ8Xo
Snf+7sqT7s0QK0bI/xc2a89VMWuKffBpA76Kv6fN3PauMfQ+aMFbvOp7f7gL6Go+
qXbZqvITS39IHXoaqAs0JsSQCFrh/3BnSi1mmECelg0+7yI4sO393O1RVYZAci9l
MOEoxGxgodDv2xXcxp4LdDW4malExCjcbI7gKhW2IuChGICeM6B368wdnbGoK7KM
yy/mbKizsGjrpiTtSYuwBiUUs1siBiTIXAd54wkBpv6xDY6riJvGK3qIWAQGDDdP
HPGFptEukzzHvB3CkaEvY0kNmhRGvbH03qZP1qDgUyff5WaJ5S651kvJyqbMFM6X
7xNJRXLzaSitNa7qtiUPm4rXVfhotIkgCJHlrSr1uyMz1K2c/dJXiJoNP5+ej2qq
+ujyUnvF/Q1kJ6bDZkq7QJIseH6mes8AW+0oopnx1M2XqBwS4VyotxyMkUV8Q5cv
jM745AYDOe+hoqI8n3wL+s0eZfiBkKLWaw/f++lo1aoq9uB7UAC/xwBeCrkRaYdO
7mjiIkTzegpaqhwzjx9I9n/j+PSky9QZMO+liERwPG3GyPL+uM79X1iOO7stiWMe
3IJc4raRK5srYnjBiB16pt6mv4+fFa/vnrikPXzXvtycqn7N2oFMxFDrTtAjMlA4
YCIxYkdznE/e3Aoi99ItDmjEk5EHjwP5DaaM69wmWTqtoQrOQuvKdgauMGiyHaCe
xlNn90PiWHutwoRLWblU+lSsnIrciVAoFfVC6T1eQPWam3HAsplt6NFkTpFkTDFI
njvgt2nHaloi8Rs0AucTQFC7VuDCkA2V15BmJN25OLOX7o1GhJa/BogxDVdoYZTl
PZKEp4Y/y6IJ7wkHKCXGsbOeGq0Y464JAOnYwUrKkKtEJQ6EEtVCa34RtKjdR1+9
sdbiqaJRbizVlvBfw+im+FHe0OW2e1reeZZIWtd7pbJoS07EJRkUQ1oYOQCZoPMI
Qeywv53OuulKQgxXERV1fLLRVTKGui2WjAqtTfBgEZ8eZmH9bo+3jibkHRCATLuE
KPh4Fy5dYW5yk5c1GfafHsJHlQExsYftbjTCBWF8UtWL47j5VO//gaKHJxcoiqsd
tHyre9zG6apL+lQEpoMOdUz4vzzboFmLDUQZnRG2qtvv1NAvfbvma2FvQuDEtdgp
cXIP22V8hfrBDj5wAwTWlm5QV/UZlNTP02UQCjmSeDA+4rKrPJdbEuCTMSyQqINR
sslcNnRNn/Kk7Wbnxo5AQNsI3j6NOT1wUU7Wdc+0cdAL51vwQy6KGNxPedWSwu9Z
HERqM/TRG8glRYWDVqzp2yYbDteuaalwKqrYh9oVWxaSLX6fp5tPA0Rw3bR95VZt
e4FQ35sRU5qcI9HTLGv7Gq9Oha0JkRpSeDcZHwUF6MIA5wGR01aLG1ykgo45F8Ai
mlYUTrVlKCoDYeZXC2iBhW6XJXzCYX40uWKVgnA1oBVT+DpuNk/M5hUADwLoc04u
TXDCTPvGFnDfVSGlLcvtATg21aT8qyjRDmKxI+DMsJEAifoLTKJdS+6e8Cbriqlk
oFaW/CgQl7slA9fGGEMBGYa9uMNWOAtSf1i4/2/04R85ZKK13vouC04biYCuogSY
XQLRt61H1crJoBH8xCKGybZGgnvrZxzrMQ9EPJ1F11IbGmSx7rHVrk83nYXvG21Q
8cydtAyYsDdSFLAIqfBfNwBGV5rypGfdchxmmhUTQMqQeJZZN8Oes9XrrFUVFRTZ
1W2jcoNzl5OKwtgKmARIdWcfvlKs8uWTzNGdr4CUmRETBstt6lDbdzgBQWzU4cHW
AGN+rbxOXOnLIdZcl9V9c7YkLQ6sv+7SmZ/FDcxCUYUC7soSZY2TX1DUKNjdfhAg
6fh0OTZ7M7hgRhPbTL9HTv2554bV3xMBoxQwmfAL8NaOztsaeypWGnB1YcNjf54q
hTNF8v1iX9MpxDPFw2CLISp2HYS/nsEcctufyjWwDo81364+2nm6K08qV9C01lAU
caOdLnhOpVXUr/4kSe+l3WH/fJS8lNdyEXGpt8s/kScai3V76ojjwTujc68JS55F
qKu0o8npKYd/7OS81f+LAY+NmC3DsnWRqzB1uzpLVdftlCDzjvhCcoHIx6dTZgbB
D+OQjYQQhZ8WAOKlf4So/NMmkN17YhGM3wAvYvUfF3PwtISI8vd08zpt+arTQLBg
5vYRGvSKGcjVlr3W/OvxdlBMttTMysLOWj6vH6fxl5NIVeL1RMYoq7NVFhpK3f7p
F5iwP3c3is7UqDMyF6aCVaO1+vauS3Wm2w6L6lBF2a4ahIqkyYfpbb5N7A34V6bk
hZO/rJOtDaE5v4QNgMnFR45EoYlqLuoz+DNRSVeZ1gkeoHXvbcy8WTubXIWu1IU9
8rvE4cKJ92HQKxwr/JQzYJUVQRGK1DA3gO7TIQi6Pv81TfgJRzBnt4c+ZNo5FfPP
N1pJglIlXut2xpBOud4cZSzKBYrVTdPJLEW+chZqP6zphQU0RMH72ylKUK32KN6Y
W8ANBCWjzOhw/odd6oAGvSH1mFmqY8I029zv6pShB/AbLUHMyq2SSHFgDTiG29DI
swYNFv25F0Q34sSTw+t4fFGur3hhmYualxjMMasr/HDbp5Rw+RI5o5w2da8QCEiN
K4ZLicyuFVE91KfGRz5/Jf+6lGanU6ojOL8k8FBYkzMuLOuV4tNCBhF/4viNK6Fr
85gP7+s3N8/6o2OuHeTI7hnA6GpU4x1GxJYrbVn119CxjqoVlSUt/FxL6IctCxZA
pTEBjUlFz5tEqdMidBFBvQ61pGpt5QTHqtjvjmX5QeAO+EAR9i9Ao8RzxKw+bokO
20pQ4YPt22fBwpOeQTU4OnKp13bTCtrHmy3HCN0mBHm99P+NJ644Sz0M6ve3rWlH
5LJagrB/8B9mvy5yU8zG+XEWUw0h3PYhaCLAxWohqCQFWKCXXaBn1lXawuWcChZ4
bPScok/+F94mM1n0WtDCeEvCCsYJ8Qy0K04R0JojZDW0xQ7xs6G32vNmEcEbW3cV
0CEUFmfcMGIIqizlEUqSng/g12hVnmYJKe6SMwLdc0qReiMJ6jeJcrxKhHrk8BpS
OSXyP9t79CBq+LUyt53FCWQ1rCzvQUnueI+j92GjGD2ChHid61FkPhh04UTQm0zZ
ERBwf3aPfrnR8PEV1bCTuYEOic7zpUVYitwovVJrsFSISziaYHncvBomXjX7cFjB
glCJD5tEXD7VKNwODQUaPO0rj3ChBKLVTLq5Rq17d9SjzYG0Tj58EdQWexTRIT6P
qTf8BIcdZWqGpkQ4VBnwbVx2rG4dMbhf1HgElepo6suEsy5kYVh48I/VIqj2Vk+T
AZu7HCDzy3ear5/0GWO4JAtc73oD36OyXGklQrRtUIuweHO+lLv9fRIF6tGipq0Q
lhKfBM2aKX6t6XYNrdbro5/BX0a7kyoQW+Lxcp6mxqFd+qCkM8pJg/pMo9aU3jKO
52r9J5m6HlYeDaLRg0OpI4CmWlBGKOSh2rEoG05YKYDqpXxI1dzmw9rJp1gcHonM
QqbXIt2t1Lp3YfhYZMh+DQXBgLTm6BHK4lWnp89LdyxXu5c/tAI2NBSc7jH5KljH
MQpb36H2Eo0w5rY15mWOuRjFB4hHS2RfmuRakaBjwsrou0T7vynOktvl868/ol54
60VXPIbReeRnTWaYRByxW6CQhyo9yNRJs+RhNYuZQHXQaOawjNeVjSP7xkD7Z2AQ
CnTgSmSFa5LbMf+Xs4UYBxtUM8Iuky2fNpyHmzVqdhCxYCGRthJLGFLSpCN6UHfX
8pNpwhJJLQCwMGbGvOAYsn7YT2b/CG1UHb/qm/eq5uRO09RqqEVvFUOTuF9XFJCU
bkpK/sMNOtls9qfLAuGC0Hl+uB/6RIiHva8tHDHTs0quslIHMbNDbydBtTw3PcdI
NT5cWyBP+NITHtng97UpGd/ov8pQfZ9PVxIQwW/zx54tcRUAQqm31TrLVyxYOhZF
ECiRV1f21XzEwBIvNMi9YjyWmoGMcaUMTTotaPue06mVP2lqxrX0cvyNEiaC19Ou
VmM9Q7zWCvAvbb8snhbg18VgBZFPls1fOGQTd56rWvXhrgDXfWCEmix38BoF5KNB

//pragma protect end_data_block
//pragma protect digest_block
fe5jhs8VDcqd3Bb7VjBcOKqlmBg=
//pragma protect end_digest_block
//pragma protect end_protected
