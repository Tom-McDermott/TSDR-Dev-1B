// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
gFIHw0zUDJJ0Rk5EpvFp1CwZOk8kC97PBBETFEuNWnn0uaNnoAbBaUkIdBwPF4Yv
iu57UCasanquicHIvKNj4YhdVa+Cv8Jrh0wPLFEkDmahy54y5z1Z8boaillM09JO
X6u/FlgHQpXXQh0/i3LSqjfWcb5RIGBWakBf2bz155cPnWstGxwWkg==
//pragma protect end_key_block
//pragma protect digest_block
Px68JAA+1hRx6lpAdIwEBWApcgU=
//pragma protect end_digest_block
//pragma protect data_block
6w5d4TCyh6TPBX9/OYFlF9f6R50jrmD3bvUhBP2q1DpyhsJx2e1erzVX7zF1MHFZ
vtu7ZWlvEexDroHXQxRRb0RsWRKDh7mBzfcHEqmpSjmaCTkeZaWkbt20qSOdCcHa
y+P9+pxcNsOFzWNzJUvjBzd1QlZJBltoHTZ9d/hmDQOGolkoh45oQOjT7uo+N4A8
RxUpCytxH+CChYzZ6qO/O96e9X19oEGAZwIGnS2fyWghT/uCKKB4JN+hMu0fpDfg
v2vzBttoHs+CyZ9KLJO2LjJGLGSuy6SD+q8QTlXqomWASymc8go8XtmQdjiw6qWs
X6KVfZPfp9QpcMDEXzCnpmegN4q7PWoOfDw1wtRyYQJaYW7sCQSONAgBJKkyj+2b
QdoaXpPycjUTZlTY9qQxuWpoiC1S8YcjpOF3aGAxxH/cQ43lap5wH07IXcXSCFmR
xsDDfCvWwFVlosTsJ6qzDUQ8o0SAWNFD2r9P+QmB4sS5gT+ImdIMp8yKkI8M0pu/
FZq5A8gY8LBbj6Idi1n6RIuRU93dbycMUz7NiHgEYmxmupqm8YJnSuFNUvBp3iIS
8qpWZ7EOqKQ7Kw06FbaMn/fvK4ZwxRSQywfU0N0LIr0ThO8VnT067veesr8XPRmL
JFqguyQVDCwe09FV+N1px196Nc0hgVLtM5qfMEVT0O9A2qqXp6M8vFv4oEzxrzMj
mdDRhk5G5UEPL9fHwaDCknmUqqakYNDwZRH8tI/zhKiAmaWBJpz89Gjl3rIZA15G
qRNyMX+Ue3tqmj0ZdV9pTaxwXL4TPTnsfNu7O/BIiKapY5I1i/VWCYbV1+SiPk41
BqlJ479IZd+OiOcJL1hDxA3y9qvjTup0FVakQfjflumZdESxa4uSzXsy3zyS7+l5
xnaKECqbeOokXi0J5oVoydRRom0l3o0DpXtRnuP8CZ4LN3tIH+g6yCKRbENsZ6eR
3N85Hen1C8ftX+FuWVB2iVd7Ks/4hfKJ2hZlfIZyxUkJN3pMJZA3dRNLdbIBpA7p
L8la3XZGuva/+I37g4wLroV/wqpmdeN+UOAHdMt2HSKPmE21FLETu/E769wjkSjv
F7clOdVzlSEO5RG6PTt8aR5QoEoiXEtFLbbw4Iq/tzlPjPqKi2syiAcmTGC7DlYt
h7jKasB16WSiIN5SO1OBrBmRom1OVC+hVMDGzLJg+EtIEZPLF//L31Taf/iEYa54
0aM90D8u9PmzUacI9IetgVvYI+Kc5Jrq/BWbmeIV7bMR7c6vHk3nCnWLQF3fzBYk
DWJN1NgIIv1MZ8lWrRoivZuGV9HR5nVSrhgYIUM/CExDytFwJtwlJC+1Uh+U08en
rmpSexwB15fhBGPNmF1CLzrnV50kVjK2TKfSlTfcFdtWafxFmb5M6y7+mWfZGNm/
ThHWnxHu9dvRp1yKACDmNZQRKN1i3BTv26iHh1qDHgC4dkqD5QrkywOQxLJwwm4d
pOfTv5kifwI9rMRjvUn0JmfSpGCGq6d4PEgn3QZLrZRoZlh3i64XXiu8nLUURjq6
BxRtViK4OimJ43ieOQIk0l5m/UjaghZ5sjBzCRk+xzER2bqOgyyWBAlJMYEH++83
Qn/xCC9yvc1hQKTHdk8jPeiQUAaAes6DUKWkKWJL4gSGnauT6awBrChNBJtFDKVH
XvbDDjNij3+vU2fuKQ+4MY5BfOAr+eFvzAXs+r9LS4Mv1zOE3BYBVqgk3vIEgcYw
f+1RDACdYdnQc/FIpSA3my/dOgJe8cwM977OLNZCC3Fd/ETQMyHnNCft1lPH0w4F
KBgBnLG7hsaMiL4GsuM6+49hZ0BIPij3adAd310Ud16PSDlEmKELwvSWt04jeITM
VtPmm52pLRaAkdyRpRVvHQgcZulUb+gJE2zFQHKyXirjEetp6tlEjXqd4sI7UxaT
pq+VdpJjz+4EapaSNOQGNbT3NUHcvI7IKlaD+60xVUUCDYL1ZBLZCYCBsdV5srZo
qJF4KgzI1TMFxBD+VD16ZfhtCmDOCK7yVJkLsaZs1ZlSypmVYXps03PCm1fq+oPU
4E9CXeF1WxPi8mq9pZ5+wZ2PtvbHzo+bOOcGaHCClccso/VKdPlSdp485VvJjrcv
N6FB9Yn2eL5MvwP6PS+gxEKHaZlXFaxgJxaQZPxZUaydoImlJKA+hs4y11GOl4to
g/4IswbFfldaUzu+ieyKr0fFEXn1ns0J9oCumjaZSSY9qYfR+b2txIYfFpiONv1v
+7FQZ5x/lMJZObmz+2E18HsOSt7Ci8vqlzB/0zepSdD+nvvDjkyNR/dnQM1p1FqV
wKBTSuTzl08/2JlLVWwX8KhfFNtapqUIKEfha6alh1QXhpKKXAO33XPwbMtJRnKf
7DJMCxG58W515spE64oB+NIrwImfX66nlQ4WFC1AKjPcZXMARoIv2nMMtkFTxQXf
weVOcaVNmZ2PU+YrXAdfNUK2cOihZmwzjy3QtiZ5cuCXGMYZOys6W355rHUM6TIH
wXBpLtDsxiPXQSWWDsUSHzJBmMif4oUSZtMnRY1m1Dhjc8piioHGcPE3EgGnv0BD
Kpqsx3qvAb25k0vw15IEZ9Ru7SAv20AF7KZG24TnvNiaYptecKMfs37s8lZ4bA2V
wUqm13D1/roaAwi+XX1QXljcMI29iasiVmOUA/9aqOgaHvdFS5zO+csYPD1J+qDh
GAMLGDWclmdvV6jnNgioCXI2ZniCwFGCSlfLC+/LIuZkb5yyH4Zqnr3jPLroTxeU
eSdy6BGx+rSAvMhL8mu/kN45vNi9eft36LIdUEnrJCmc1XRedoxtJfTbRkT6cKDQ
P0FSFtaI6RpNI454yBMszJwJf+na5pfXYe5yVFjguxaCDB9cPmtbALJV0fBqB7Uy
ovYOxaLF6enC9nDBit6GoJZ5TZhosSOLzZHPGTqZ7QuhXe31KZI7cB8VrOGiKW+Y
QyrCvAqedMixHy9meTSdyUuQhL0ThoaXHn+j7toSHiUOP7kjrg//SDjzXJrEP9D/
dwKuxQ3s9eegdo+fEzl4wC5aN5vwkC6RfGkR3OX2y3OJSSGFiU56gMDHjDGivULb
cf66ZAzJYIGM6ozUPyz4ZkT9WZcIts10BvoL7440/eCdMDmfD1fygRYGV8mXsujT
0yhdFEAr7PAxXkPT8JzcNj7utfuPLENl7U7tYFEmeby7SziQAplglqTM0p9LtkPG
J7JZ8gttbgWIYWLBmYFIn1hzW6fgO/pe1paAtrInEazKDvsVUYFSrq+GbFA06Frp
FHGSBMTwrCOPQozqDG88/zX3FZTHC8wRVCsWod2beMC07P4r2ZV+uF0WcsKLq8AT
WC2QEhkHPEO28rVsjyfg4waVVDafEfSXQFBde+7Q6byC4MG6dFcB3D8SV++JWnLB
O6bA938py7MTWP6251gvou+xux5BbzzU2sopZVOIOnCcQaATDbEs6/i1a3mY9wIH
QiScPJ1ZV6ZdXTyR+TWnCkN5vY8CQEcRMcwn+MN+D8fdUcooeZpS62Hy9o1RmOzW
GtSLnDPRiMIwUf8Snv8sEeH3xiEtDihn5e0VDsRr04mFV56Q6TQ6sx3H/mn4oJ6w
ittrHgBdB/wQXKZZvG0/7+qvxW0/i41Mmg5KRhZt/hZJZAqt3Lsvw7P0qX1mRJmJ
hxE9qih2pRBFYRSehMcejM2QlPxSz1wr/32WhNKtR4qIJa+fROenb56G1452lFli
J2vQ5s7U9cX6oQl/ccjy61AARj3st7AyWjmJiEd60BmJkBTFoLrxgU4gwmlxpV2a
U8XZEKz4SVkGkC1nU2wSv2So65wGR31sjEvjxp2CzCM3j1Jj7EqT1NDcs0EeUzQz
knz7iPvDmIGdbCmsjBnGKopHoSPOiwLATmW/uMgMmm5SUqFR62qBRPKJY4toJTXe
D4OQg5wHPd8zL0yUZxWcOww0U8DzCpte4Puit8NS0IfB2wZf7PZuWSzDN6O6HZe3
5Ya5BdrNi+3eLmM3A06eeSnyEzq24FQtB3jA3Wpz7kXtKP+8z+AoSd5/7wDCSBdF
H3et8Ea+av8NvUa1/y4ACGxFW7Xu4gnHaPPX/epfU44p54HVJH5tfy1yARnYoMjH
1cB9oSlofgMwpvD70qyVY7nK0S+0vZ5SXh6Q2dkL0aLzFnsta44+mPescrkJicGE
uDMCPxMkmyuHgQBSjLSbp+1td2saXRuboc4FCqa+NdbQcTEJ/ip50XHwz88F4zJi
SZJcW+op9lB/e+jxOoa+t/1CvzXm3Y9JpAiGjISHzy3/NrZil8kh2AaFmudzuno+
gFIMROvdZPLtw55v0FV+RxNPQifsGvsmM8/F/DKs8En9mfZVw9sVC3WwpqjXnCv7
MAPyPbNIoSj0V9n/BtBSCytDuYWd8CZe4yByI/px+JSP1KMn4SGgCBrSy6O2vUR/
+MRBFAlF746Vs00Ms08p/A9yMCjemnNkz23k62wyz9IlgzfXR/NdtXfqlhAJAq8a
miZgy66ccTHJrobVsmUlR+cLQ/RpyxofUuNtC3SgERFAV1wz1zDk1dqKYIJq7wgy
Q9bILeduUbJ91THvqjMdkMlhj4eDprIjn+WQt+eq2JN0HY4WCf4WnRX/99kg9oQP
iMpIPEoYGyG9y5hUeCOL/omf+WWQyEh2iAu6/eM3EhgIusb1kSJIamwvis/6IeHR
eC4m7SQssAfkX8xa73He1Ytj4N9SYYmyMl+af6SAt2wbV2UuHEpFqBSsu4TMEYoc
rASjgCQ3jpWRJWy4ORnAyTEr/ZaBK9mERq2CffFI01Z1vkQIo12DLMczfX6o4WKO
F8ZHUMSP0wmz5ekjHbzVcWeP7BIkPVFNl4dvenHB3kM1qDVghEZkkzvviBR0SnFq
DrnjXGm293PcANjMPRJCmcijTT0pDo3Pq0c44DnXIeHIcxxzXPujj/PjhJmCyGXU
pEfZsoINAdQLpithMyrhjN6b9E8f31tmjR/WDcq565718iUHF0x8tEtHWTQQVQEN
bORKg/Usn8hMxuR+PK1yDPAAOjxcmlwv9Dneubye/PIpZF9NI3A0aeBy7haGmEyd
LdtDPDiQ07DVT1qGA6k0DlVEz4Am+qQV+xYKckbV5Myx8/jFmhal45vpZMP3r5ip
o9sr0/Ld2oE4JtULKTiuYM/wx/00wkm9/3IsMPaeRhJ18KZIO3dNWoKwkBx3KDUf
uuKCD0zf/7YUsPW9jwZasBXxybX324BSgbBBwlOC3DXqwGH3yyN8PRLqOKQP3YSb
6x0tQrR66U89gvUi+jKoaFrj1J8Gwvb9LB7wIf4D5N5+RrdH8ASG+tBPm7Dj0pdO
dYNZu2kuwE10Bdfv7lF3rMROMX8HCWzbo7xTkjoPQiv3n/Xp+c8FyUHduL4jeDCr
Amg5Xz2lnljdpDCrRQAdR0/K7svpNEGvY4On/iogLyZ0NXeDMU2FvkRWKEmHzIJ4
//V3B3wV8dVSErYTfC/8kHu1Gyk5ASZjSzvucIfjIT/oMAbBiiJAay4izNChGPp8
KMOCjyCtorX6JNhNwyJskWgbws71872fUBvt0gz7cDHplO9UHHn3R0NHVpcBwdSJ
Pza6CAuUiobf9QLOs3BZMhI/2myxfMQ9tKBYFIQo4GS9Z5+EFIhDqqQnx2jipmuP
PRVdlYiW6kGyTeKajylRplntWEomGE4Nyx3Wmbncgivp5zoxLHHGvTX0akIZzt9J
Unu7Qx1KFLvLPVGJ2V2Lr1Du17XPXOJwX5oz4b098WXgx8FbIozpNTJSKijuMyLg
y14hYtP6Ar7QRUu9fGImHub8WcG2pwKUvl8QNRmRh7bWAFB9XZUm7joFiQmcmRlw
iLyNm45EBLPgOOfRdFbOFzbOigteTewUi+BV6wyCGGQeFvFq6paPAwkg28eyGRl7
IuoSohvjdp41VFD7p8r8RWPMif+993ruG7hvK4JPx1384ntSxFoc1Y3Y3ax7zcVd
ORgeqb/QXKHtWYHKQvJBKMLciS5g3Bd0aYz7mmhD9t2dSJyPFYO5wMarPEV95gp6
e9hBU4RM7giTZhob3li4CsEfNJBKIalVP8Q/IiDsm77zyPCXMt/NaDMhOn26zMck
xZGkRlCd5HS0cD/TXYJuu83oO2mciFffPSQjeSwcSy5R84PliNbrxA8JKwbNWIfW
ChTLi7j8ExGGaUJYGhP/4n+5H5K2649zqwG5DOAEd/XjCaksN0sJZ97B068JVscp
gWAtom/A5Z3MEnLzERY7AmCFnoErapopHTeIIjrUf1OQ+5oNAgRcnDc8cI62jDRN
fYyEbuZJnGI4fgIRxAgaJaPr7qW//FDEiWyW+QeXqYSxgxBQWDdyO6C1zk9sQd5O
nNsGHzjmC5Iz9OuPKOlNjhg2hZzC64G4n35FlQ+PQbwD1578akWWYk8CikwJC6WZ
v0VRZK2H+1dRC+vGm+WraHzuceDLzW5F3Hh8IXjITL/8czuBz3g2C0r5FHhHZQ7Y
7yGfHaoDGofeTaTsTTp5eqqGrVDACTYrmjCtleeFZFGCHpWfu+oK2/Z8CzPl4uOl
LyRsrvhf+wT0VmKTqsn9qwbH1LVyTEttunMseJCFHqlC7oa481cZjT7HcZ+bJNgU
ClLUMCa0V1w3w7aMMwGkmaEy6uV+WWHTmJAFJYOOM1PvGew3xZ8WxCGURAYMuf3l
enudjS08fDQ3yVGvq0lldS1hbpyNZZuG0POwNDG+gDQKtrVQ4MuychSbhHNhV+g6
NAqF0mHo+cdZE5xBAFP9bRf2H1zVDXXvDkGvhvtg9T6FXyOoYjx5NXyJf+kzUA3A
mkHmnyzzOGHdclwOcvAJJ8YR+iDrcviuWq8RldkhjzegT/BdIwdtES+I6wvwjTy3
UNO1VLONP4+AoGB7MSo0KcTdm7oNdCYZD/+dcYqX2s0N328sdMorAjtjKMrXrrxK
eF+zCSXJaDompLu5jyOnza0tHy3nUNnNPX1OtbG9aUTs3WVwieZO34anSgfBQrLF
0SyXqZRxeXkbdREk5B6jK7KjjgBfmr9sxMn8eo6l6fxtksY7d+HFkDzI27rxrgnB
TUObrj6tbq8DYlJ4pi/TnIsMgOb62Bsae8DrAQA6n5xaWzqSeRFfLX87BdKWN5qk
3Bg6IxZ1uDTn3NaYYnBSOelsJ3pknezNLWtNsZcMyhvnRepJPNZg/BTKydUsHkRB
5x7UpbcrHjs9s4hcs7Zt1fhpevpAzCJX5qSC1eouFctho4Is9a2J87f9wzuYBHQt
MickrB3zmoOzn9gcTgQBDmx+2ypQCgS8qQUIWFd29cbxSNUz5WGD5Hz3i9JJYYvR
DVMiIvFuSfCP96JRYRoj9ZuRSOKbCzPbk7D5xA3lHUHqPk4nqnJT53sFkD6EbABQ
hXsz3FOklyJYYnHnf1VhFUE4gjVkPNt2Q4O3gtMsH2XWqs8zzMGUFssoiE0ZzIj9
iGyFZv7o5zfvoa2kr5I6X9LBKGLGTtsTdb2h4PX9VBQzJU6rcOQK9JUpxaSyB6rj
Euv9c8q14oLXzOIuF/zaAd8Rw6K4IYYb48rwUpPTALREsKqlSL46UNbd5tQsnJNI
jCxoG3eHF72uNSagWhReZ0IIZAYAGQJKsvEKolj6n/H0o4wSdpRulGuVuhu34lD1
s8TSQkQBjxnFU0+kF3pRor/ok1fAtuxxWtYBFZzucEeRMmyxDIAcMoZ4BUssi55N
ae4cLMvq30ICP6Ox5Phb1QZOUvRFOEhEhSzH0wBkrwKXQrBEDG11KhU6qnbpTIUV
MW83c40uZ4ExmGBdWHybUwyiRuHxC1P0CaK7pMffWTLqtYX+WQPHZIN80RP264jj
3gadzsOB6ChWMR6WkfpzKu65JKk5yY8kfJVpA4f/iooyEB+SLpajEOv9IqOXg87C
GkVpk7xwwbroZx1WPsJ0dllce/WUK3ZMz/Vl6nzF0dzB05BGI8UEQkLoJh5VSeKn
TTJMY0JXN4LZW/ueAgC1xIu9LNjXvnesEYoCfVEqyoWeuKlxxm4s9edHV+poZFZU
8StACbghraTChPsK4PeUkrdrLneeocjUS+MEHk+XJWMAWtXQfcSXUHyuO2/n5/RV
6J887vvF21xVbfbQ3OAUbV+J3iD0zBP48achRQN2h9q1rlFqdfc4HdaNwWz8T/fp
VGc8H7ibt/hF6fVcwMDrPBnFuzDUIjU2u0szhJ/UZhozqyKQcFJ5rv8A1HbNQzHX
3zr6vv68njdxdI0x0T+b/wkTPNyaxiia9STW4FT5jBSEVHqGmoUCHu6mQVbNTEH8
8irsV0QAsm3ZPkrvstnzT7AF5rSgEFrAEuMMuY7u7G3MEhpFu+vzNJTSCsl4H3q2
O2FYCMYTXPne+iaGWIfQGMuMUCZzr1WplM4U2eeJi04M2M27iKQJG1gzts/Tdmvn
jwr+Ti8PZTlHn1LlGSy5vQE0tHJFgh7nfAqqw8WmO/O/Z7ruS3lYPAaOQNoGnYLI
jJfEgZzar3Zb8neMyLCUkuW1bUzdBoN5Uvv+qRVDAOAXH6C3ewz7ESlug8t9GU7M
/+VHweZlM9r96mZ4hkVbHTL+fCt6JUguOw2DRtFvdYIesJRHC+Nci4DH5P5+YejI
KoX9OOVDh67xAWfnz/0hMvm4L0SUiWGe/e+qpbEJN/xgphjJUkEl3jU7cdk8kNgo
7oiTDoaPdV2YvLg9u536hzlejTVM0ARVPAq4s+lzO3ybLn9zyeSLTm4dnY5lfXAk
sGvuBgKoLv5QTA6zanjVrom+0CEdiHRmqlhAYklS+0sZbouXP0v5G6RHNQNVgS9E
1jM5SjUulKG/QKd8ttRQs1JIf7WYcALf6fya7E1eS3I=
//pragma protect end_data_block
//pragma protect digest_block
HbJIw6GoGNuy+BJ2faWS6nfuGnI=
//pragma protect end_digest_block
//pragma protect end_protected
