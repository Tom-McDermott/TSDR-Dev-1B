//__ACDS_USER_COMMENT__ (C) 2001-2020 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
//__ACDS_USER_COMMENT__ ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Jmdt3dE1+/+frnbUGdtDTiDyXvIZ9/i0po+bLdR26oiEMHQQcSPgqXl0Kw+vY0NnR8lE0G8JcCOZ
dqzjX+KsfWv3KE2S6J9AtmJYI1obU+hUrYc5xqt2ZJNi4XVHzV1njFnTNBSSos9AX69Pr2hngxLY
GHF5TEjAnl4fFixgl0Qc8V7ClWtF1AuIr2x8m280/7Wj2MSOuk4146gLOK0k5GHJwHdr1K73Bfk3
qMLYp8GA+ASIZy/HuevHGgkKFuv8I/EcC/3ChItnCtJi0nZ+4DinE46K962dSN2V0bARcq1IX47l
Y2/uYDH3uDPrmU78BORLwB2vaPsyUqjOS9Sc7w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 12256)
SMHJPRSRESIcLg0l5rbJADCnXlJQfLpRWizCb4lAGEP46V0modCoNHRUcDfMkmmnKOPFvBvtWRa3
j1jH+bteu1I0mgTndm4GbPncG7CbOmm8PSn18fQcHfAHcTPdaTK1d9IsZlYvyx0HOnMT/hGHT5w2
qr6kyzk9vtOQTouJlBk/p0FKVC8EHQUhrzct4G9WDXdCKGXJwTPs4SeJ23JgN7EbbklFbtC1pLTF
ZTsq8zV+4vkSpptQbNHfJmMW/2wc2hqY0bueoeVwhc6qUxQPKgqXfq2ktQ14hwKyiZVK1Z2BB1b+
jCbiZIpZv4Z+cBL9uK+A8/099+XoyvNzYH5GTL5/EmA0oIgifTMQNy7X9/tDrJjas3DRvtYygEEy
e/up86wsudd4ZU6TaE0I7tkdrjQTIy6lvIMiTIoyfVNpMbIF7HvKZP9wQ092rWOArjs+O9i2ujN9
mze+CtuLdQFhn7zgsVgxWjjqzQE+u64iFLzEsTvFaKQ5o+nGrxYEf+zMOfFGcFQLK7xznEUH9P/J
Q+sCAFxqKp1O/Ak7Zl8XRJDmoAUGjnvduLxV1oxm3vatxojgnSfiUnQ5UwGW6xfjrnIfhQb0eAaA
XfXhl7K5nYGVsRo4ANScaOLO9p33fqOp5xKRHxXuUzw9pL4M/+UXvXh1qCrMw/4c8+mp3QkgPj+M
sslCs/URgCozRVSl+4IX/qmsUjrtVhFQ/5cPvRxYhFz9ylWNTU6peV2NDRsq/bUnZWRHxoNasLZt
efbDcOjts42o2acLvd4G5qc5k82xyEb/OrG7VhoOjdcImq93wPz69UOAeKyLWAksoJR4zMSyUp7Z
nGk6JJZEPD1J8XsKXET/2fu4jYNUXFJa7u4g2HjkD4suKiXizEdGsMj85OwSO+UdM6axxrI/oPoa
Buqgj/NmMXKfQ5EMxnZpq0cn5ASr9Vq1jBo540hfjWnY0q0z6CMm0/loukmk33vMEUFbuKcJkfmN
tiulrjYwRK24IA2PrF9LuyBLiG3kuV7mNzg2X2TDYK9CBUOWNO3VH0NeZWL8NIZsBmwwOiA4hsBm
pKmarnSj0FtU7Ntxqo5cfzejEmLih87xIqVGCofZAoFToY4WRk4954DlZ3Ew0zFXzIg7likrmB5A
YnZpzeiART6f4M16kevlH/nXnAiQQTDkvZPpWH8I2TkLj3Wll91Rz5rRqg9oe2930eDYMy8p3Pel
dLPhFDpMUOVrU0OPlouViWyqilks/ghQ/n9nqsTTOTd2/17TPy44abU7DdRGxUwxsPqtaPO34Y61
P7AoaJ5bQ1/TQUp3LxHSXRuUU++3KnzShbgzV9kSYEjLCn3qlO6v4ACzyOTK8l1nUzUziFkbzJXs
30OUGHN8k1PPfEDkTgXCZRa1SXfXNAdDQtIgQOPVlA/o3qS2EMsELg4J31yJmCZQcdXXhW4VU3I5
blDRmjpypzSmj0OZJZhIpK+0jqBp6NadYVf/4GU10fAHC5Pc7DQEg8mUmpyvXB3rFlu2fSRLUNAg
MlV/PokLufbJJ0ObOKqKByS4NzqZK9NV1C4HpEF08jiyhzI+Jj0FpCM9zgQItqNZCRPaPHNZ/jSQ
bYhHgGRwz9Cc/gVU6Xb5QlWOM2yWMyPQg8yegIalFlPzfV1CJsJ1PD7s1Nom3fY92psVok+7YTCt
vltvu/JcDpr/ahYceimjn4glHIhml4xC1u5/HMos98x3ys7ZWMlt5A8Yq0z/FtznmlG5dcv0noC9
2soe1wscSoDUaIF8EgKwxB5B/X7e/u8Rxa1IcpJrtWKgOoE0JBRCs5SDCvu0PZ1jbn2aLfo0tz2e
mZvPGC/X8JFkb9nQGe2GH56xnu+ZuMVWffjv/wK8XmIRAGKFEIm7z0G+pdgk++PeR2epEmTrPsvS
7FX7p+7FxSyHnK2R5orRraizOchIk6wzryx3aTa/Ah5IHDdwql2fkojJ8IMGIBOxkB4sFfiApPVK
TYYKV79WJLzEU2o7fe4GArMJQ8AOssn8HHAc/Ql15h5kEceJV0McgK6VRDmazafoJCun9i5oZPiX
yTNEpDifVYj/7LpPYlmDby/qHTaJGCQyPBzeLQkmHo9giMHJ7z6sBb3j6NE0nTFz8N1+gTBrEQFD
ss+D8XHGds7a5IbodnkAaiC4TT+4egsXbzoGvI996LYlKzbL1JEptPAs6gDlo9MYsW+PisC8a08N
KWMc1enY+zU3R7G54+OHzk4bj6N0SruKmu10AmWV97YnyESCIignY00HEfaBF89gOfiCPdnAFmJq
lWlI/L2+TFWrnk8WVQB9LPhQr9TlO+M4HX2IeaJ838dL3RSof8G5IijavFDUq/WEEoOmdgLbqKgI
mmFc6aFH+AJFXTc8Az+RhHmENFfIUkjvCOE6zscdbOCvd/oWaOVRpwmQK/uUS+0CCELgO6pH6yhV
LgHWzzG8w+gFemR1+Vn2/Sl6h/SVniNhK8GoxmsWier4BXN2H2Z7/z5yeLEwwDilX2aibB6aDMGE
OIYQka4fjFb3xQNf9rvTYkESvWXxhqkTxVMV9mXHJkOiAbfM0/vKQ73slvk+YBSUFH0BfnIuZ0Ib
w50i5C0O/1vQv2lDQH5U9rm5IiH81HV56DWMyK0yJXGe3cuZNA9EqaFXXb/fyv0KUxWdW4UqoFtu
p3wzN6YemTavtssE4axIqINu27yVVcMtg/ynbm3o6fXx2S1X3R0E5AMhT1Z8BS1d76xwNoakyoMv
DjSL/qKL2F9ZwKqoB3DxX7KoXltKhqdvITHL12RkdQN3Onjm5DpA38k2W64GhfAf3GkYFXIYFoBA
eAlFA7Q9pn0x4fgFImBQsoBYFYc6Fp2NPKqfI8EAsJAbB4ks9puw2/Ew6oeuu0YkQV7Xx9a9rSYe
oLTLmmK7wxj0cRZv5lVcqu58bP2JqZWVCka2hrihXlhtdZVw+iA97GUntoxXCXycPPuCeqa02au4
Gf35UTA4FzB1vvk38HkO9D82JRLclNhjhVncrt9t+0tasw3+R8CNG0mgFMEL8EhEvxvYRt+LVi4E
ZgP+G2earSobkw6OBDSjJuoLWdQEv9Vo5Egjh3i7Xidk6VjoEo1mcxxGWMOC0qe07d6H8tF4yxTo
wfXVcOh4L/Vg8J3gOoDJALbqCEl0kmKl9FOI5V2WL17bfdb9e0dWr3YeQYqotjREKOgjLCedz0xT
RWgHnpOKLK0CUakClEVn/flGwAdCXq4/kKcOQs9NaTf4+xk7SsIIRgiFYd0w2HGbpMBwLjMfF0EI
T0ZhFRP0YLaVky3pYVt1c0OVOJ6jTHoJYWD17PmmosgHnfBLctf557JLyIFQ1yd1RsvjbBaMXI67
e1/pnR+1O2lcHMUGg2sEcne83OH2Ewosw9vp9dE+J/7cr1UcdOV2EodKfFBzJucHS2bddsz3vQKe
K9PfRpf8ogzuTA0co3obwlEfh2p6jAhvLkVc9d9ShdP2+J6Hu4oxkVoRJ03ToGnpvUQt/57AK+ib
c0BIMkon9paS1aNPv+ZrLQezsMgD0YL21FY26WRYrh+hjkqJDiXTr42+Jmx5TQ6MIlJ3G8jtvfCb
1ss/V00ldaE3kifRgGv34Fcehhj5oypXhWwqN64AKTsfBdRRasinQZd4mCih/SQaGnDDY59mTcTH
8QesedIaHXBKzUXYlIN9s4XxmHyuQx67JuvXvj/Y1vbn57RTE8DVSe9MuJjT938HklwpEPAwZxL4
SXOFc7KgmeeywhUYc81Lb4+DVD3W7gkZrLCa8HIs99e2QYRAR5eBKyV75fiJevQYOslGFCCyZylJ
tZGlBXHKG2RWeACQhWRIdK8SBUpESdBkmedMkfcsVi87wh/sc588oL5X2c1hKgkLLI1el0/OVhDv
YheFWlKXVFN6j5lE1/UvUTDNqbp/FudGtxDh4gUsKn59gtE2pgQsDk3mYmB7LRlksgSVj3K23yyQ
dDNCsodAL5xs7FHMmcFc6tA1zr99hkGoE6VrtHLWvxDf9Bo2jNwfb674Km6Rl2n8nhe6+WolPYFQ
UKaQZMeSo/3Qkxxa4HhHMMvGFUbCmVZM5DQNzjsMmYQX/h9o7jHpkgrvM3Un167bzhv1exHqVEso
Lix3yjvc8vi8aa5cbGj9Qy5s0AGe4w3BR/FmbdV4XvIhsFE+wHv5ReD+jAIXtlFH6rk9E3TD22YF
g7n3DKXqo8jPTrPBxtHz2YcP+sMJvwTEqVmskRGhOC38GemOV46/7SbQ8LxBD6tNH/Ky4EZWx9iP
mjY/E3Zfgczvaam5smbWPBcMwwp4jvHp3wu8nCr+xzTDkXKoFUBMpZjQeqtKB17/MQ4cPU/aPiT3
7P57mGtQnmwwdasfn/C6Bee6HWwLXAuvClPILcMu7QoeZPbNi3okKylr3N4QZrJvrYC80oOi7NTi
Lrop7PvBLyONbNu76HDKdbnQvo6sfsSz397Zn4tX8G/we0/VKTZziu5E3Vmd4GwHtonziELZzo3h
2Jx8BAU9uIuJJbWpNG735Lse5ZiDb4xvxTutH+J1G/Mxo7YdK4Gkhnqa3KNFTFyX/23JATq4Kme6
RtedOfm9hqOhp2cwAegkOY5vLIkx3iDABJWi2yLmNtbzgA3s9nfrfrFqK4kxjRhGL6eMlJ7qiyw7
4110AbPZ67xFolEWiWwkatBdRvOYSXiLZodt9o/HXU9WJw0rxtOyiU4Jey5FCurbZVKihcUTu3uH
3E//JJmV2OTdHPEeyn2ZTUCdaIZFA8ekUB+lnl/p6dioY0qQBUiTypIvXWrjYj6wycJWRMPzjhvv
biETYojH5W9Rb/wwGf8a2hVjLN0eAOWhkG3DKGTWxtq+GDQwb38D2VBOqfJ2w2zU9yQR4zHd9Pwa
C9QA66IZ4heIDmI7gYjM35OUXp+LaIKD4PUnM9nQKCWRWtwzNioUbu9YCKt7KgB2+RqTczfRnft2
tlq/NKfo94DpS3TMa14A0DP15vO2k8XEMpxgqguRssv4P4paXIi3ls2W5scPtPc2XzQeksaqPL7G
E3GmGkkPNxsgS/SD6zBghFcf5haquoqF0p+4mVHUl48tWoiwn51V1aqcKH7Ie/h2JQForjwDkbyl
hzmeo6Jp7hn1xyD7ESjgW7EWOsX/6TKj88px1kNH14zEg0NtsA1lnPEpzTD8yoBt4REsoezbbtxm
F7N4HCEMiV97rEJuRMeM0uFFmZo7maDpvFx1+UdTXvp1R8ZKe5AVEBUdJAZfTjR28jAcCNwuS+zR
teirxPS4z7GbCn6UrXSsPsr8KHDZm0ySEvwVJJThWPSerF9lVhb4X1YNSLyEUdWZfEeWE+Kai2LE
h+hMFbpjHyJ1K3Ya9lakKs4RNbxLRjthl8WAEpN6Bls64DgfjbVCxs0iIbRPR55TAWdAWASRLLaj
mbAmIVS+st7TQu5B3HpEKqF7Xfabg9knjbM21mhAiobmVL5a+8sAv6saunBMHON6lVhGFph+A05h
V16qbvmb2SGtkOqbKW+DMUxtPRdS2MiWzILx7C9VgCmyNajmn6/6JBF1x8JFwMAWWz/8kN+2ldJG
OyyxZIT55Fmnsoze4/X+aD85j6AJmErq3o9O8/kdlig0oivjdzL0rXeenhbsTwwMVfiC9bnr7Dvy
OXLyt8Vbt5pwQxqZxnS7mkwEgcuSXjpcIH67Z2z2IrJRf8FsqHS80mmUFgvBdkNMWQfSKDo4g5Mj
XYEpJ/R51rvD7wR2vP26a6e+PtGo3qhaKmOJD72QJsPEBuf1DN+ZqeCiQcMdxX7qbxpA2fJZ1THg
9nDvaiAWwKPW1M8PIeA+NinmEnI4rjLNRwSw5uogZ/dB+BWK61wySJ4QJ5ZGDmDBeZuDX7F+oheK
25HszfLHDpa9m0Y3x0AM9+IAz7eC0KX6GaiI6grlJT6Lq0czld5oFfZHe0gVVvEj4lxFGNhVFiVy
2+sPS5mnK/kDQXIIfXPgVcESQjxQLzwKjYjp0zS8iISP2UzatkklS7Cn+HrAaGudyIbt6SYqGh8g
SBugMOm9tBecr4wNAgrUeacdUpicfjdrkd7gbuUaY/qEkJzTUFNt6/XwdsK0e2dyiMLYPYDx1bHO
WWHnmKLPDsGxbNI3fhFpLiR0JuH1QXtzipyz34FXIi49r5PSt4wFuE8Y51hxz15M6FBdYs5/r+NF
310M2jxHbr6wiHqDY3CFBOMwSdL1mVyHIKMaUNfsZYTxreXDSOsPYEneFjp8d+mCxit9XvIpQjwK
fp9iWHy/UiB2YyLxSc/8cyisZJdCTbVpn9d+RTLiSUDRqa47I3tRj6k9kWFCm7kIyj3PiHECjRLD
UZGCHJlfOe1ltkt5aeT5JGmDYoPFjBLZkgFJFazBZ+Zk89RVVr5UibbN3cyd5d+ahbUfx0xZs0fX
1UBl9Ivzkod9ZcvYM1vxT5t3TthlYEYA5ombnWapFp5bMJ6b44a6Xl9ZsClst6NOHcycvrOAlarc
bs1ipQ8egjW4TjMNaYcJVwoXhXsFIgRtUicA5e/DKdbJEkYV7nxkoAGGdyKCCB8jx6sVLccgtNG4
XIhoKr6EvK3QoxgiCAnvf9zRMSGjmGoD5D+EDOazysx8GkimPML7W+Xtdimb1zxKma8U+pXR2opl
/8SErvW66Xe1NO9r2vnsnI9gWwK9bbfvHS/98WvfhOpk8kEnT5DPeoQwY2/PgdiyM++6TFQPC1UV
Jhq0ZrC7oKhqBfYUiNCjOulVdKPfp8r8v8hgLWFxyDpuo2Ik9XEVGFIxLBdhEyObH5ofWDhCT1ZM
TrZlxV8fyhPzqmgepLTryXbPUVjvtcaTAISJHwxZIZAgSv549ZdrjAM6UDOAJvQZ+yOjnbH4wZ2s
6x/Kv8gmNxKa52qcNHP48hRrPAXJTvGI88IW9Di0Aq99kA6zj86dWm9Hq8O2ujLCbwcwX2Ve3+Kc
TLp+fEsTTRrd/uSSiRCEq8k85oE+Y4TY/p/pdAzTPvxvxzEUzkUq8dCLid3InVL9MkxBvPxx27vt
abAWs8iZ4Fo4BmhihhHQpN/rCXuYb6TbM8kFeVkHdyoM/IROAqBxlQmuSrLP4LeisVdQ5LPyulp1
BofDT0+kbDkSsqGNXGXck3BgVHzB1z0w7SGT2KL7NDFxY+37RpGy2LTqazoQQcQTTXY+J1BgciaA
qLrJ4cmh3XXGMllpJh2VKTCnegCGOuhTWKJ70GMWFiiavGhhEOjLmgB5bd2MK1j0Diut0Q83EzOP
UkTXgeKdLX2+J2nLTzn5jpp8xfNJYm/psH/q/x/Ot1RuLzbSt8TDqtGjcxe2F+8fB9mICqcbszhm
pm6ZZ62qnWTdA/09sYRi5R9H5BLkxl2T8bZhxT3h1FzzhGpX9TS8qkbpPJfHqZqoxS+93/ehF+br
WG55ef8l3edeujV/aPKfe+HkRXJeo2DNyPdu6MS1hsrw0sefe1nShLSdbXNUYblGcZ0kjViA8Nxg
6Y2RAboI902OiBZIabQu2VFwfzmEyZlSDd4a38JnVaGhnfGvbtrooy0dmfl3/CHC7psubYRBZnTw
BEB20Xi9XA4tIPxzB2X+9Pmaf+Ahur0RUW8mjxfLe7VAHb0wtg/vX/eY6hX4uEDt3MGtu69s2SAO
yYxCeF9PDLdJJT5E+arVsh221bV8L7fgKO2QRUtwgI0V5IXX4tUUGb+mUAT6zJZKAIpj98tcqznK
B1K0/CmOFJWnMsu66l6pyAR9HV4ygWHL3zPBkTBBZqf3m4WU2c7eVtOfwlmpeSVVsjGIX1+uoiul
S9DgDs81NPBa/pzGAebFMUBsre4y8zXdA8eG7Gb2uunpvtgwOEwWDku4qiVW4Y8aZr74dEatIhAA
K089rIePQceQKjqm6zNNSIbtMvIgnvbW4aSv5itTWIu+mQicQLw9saci1avjoh6PLODAV17jOIW8
jzCdO8uYZF1nA8XyzaBALbmn+XBdni/Nr3GlkrwDB9INhzvRdmf+dCRP1doV70dnhSyIXs8GzK2W
ohTVCjicHyYNfUurxWb07pz7NIuNaWUJnONhUn7W1Sm2qRRdinaSXBAWoXc3LhYFCb2IJ4k1UM+w
kcH/88PXbrLYavGq/P9E0BfH3Q6+dHbdsxkDTPmQPbNYEbkNBoJhJjZdAIv2H0YaPyFfx5QLrO5k
CBS+R6tz4oZZLFO5Czt9ffgfX7VL+5a+xTqbP4B8F4AXVjHKBck+pqOc8LKrTiZT1qKdqvnLrDn2
UCuRNvE4BnC52YKfJUr9sT9W32mWB/HCQXmXQ+OP1afHYxSkl/Upvnk7MEc1w3zQQXFSw4aKEiy8
x+boq5isM4XyDzwUv/YvyiTY6EujwwVU2jUHxNmUAjjl8HbLYMoBY1lsjiTOFjksKDt5e89EhInp
9VMz+vG28+IK05LsyXzxISsS3b5X7h+Mnm6OiL1zD/xF7yJAXl6Ynz3Ux5f2L2KlJr2EmvlvrYtP
7JRAOVX9kXCp4xDHbEb74bLKrH2hZGB9pJ7HoE3q7bvxxK5QgueRNClkklAyenhDrsT5//GOnvzp
lPIwoBfb5WAh4m5RJalDHxjkEw84X9KOzO3D5yryzf2TSTIGWbv5uIPwM72Uk4XqPO9DhvPkQPAU
M4e9IPfFnn92yyUrup9c6LOVYX9JR3e7YCSOOI5p0RwroSRghbFdUFcAF/U1O6BwgThV3TWUpkHr
Ju4ARmRDz1AsdlSOpN8x1jmpsEKAWt1zr6U1k9pWYeCz/W1POROKjmX7L9icCPkRvF5jJ9VEuhnW
QIHtJUOK/vmX4ATpmIcgSYX/3yOofEmOOwkYQuGgRRwU53ttUDjEj15VvZONIquYtRVbld6NIiW+
d9VnmW7L9IF08X8JPG2S9TTGil3q5ZpwgRAJ9+LrFu+4xCY3XXvuQGCcdPqBQel4MBKEzvzdVyDI
V5I5G4blhHv9vZqghi3omxF0OuRfXE8TKWqO+ar2SRIzfAA8iTPn4tx2wWGRcgeopl0u5Q6heeJ1
TBKN/hfvWG9JFTnKFB4XNibltfFWUrEz8tUzds/P26y8PCgdoEsBoDfS0IDEvNBcHMezVJCj3eSY
VwpfoVKv93llF1k3sb8xURbd1aHTQl2PdHGJ240qU3PjAh1YgcvczTBgMw6b9IipTwvOjZe84hhx
6zd1ZSg8Gi2DdgXIMME1u7rQM4wMb1jum1FdYUh8tqddwXmIJKh+5m5Z0Rb9CvNuwHsuTqkEapiF
51ocqB4HvKREDxsT4RifBWEWz3PuFBjiMrCd0bOA1JXCubSfJ51ObEJqeO1nqEWgrXTJkG8PhXfe
Ui4pWSQitensZ6DLildpspc/rXUppeGPPumEU2ByAcjwTeCIvW6sY+7m2bQ1ZA9bnqD0Y3HunzHX
F09OyJp55bRoKK7OyDnTNGC1Ir0Ncw9kZqhdoYG6fj78p/RHiL8Wg88605I5ziOicg787YgX+7P8
jVPwUyzpaPr6eWdZhnlqEoG7rhbCMWK3rxxd4mtUym5WdREk/+CHmWRgm11H+6za51bEVsIu/TBD
P02HNL5VglQNP8sLxXxqGxKLcdLw8YF9xL/HTQ5fgpEl2HFRvxBewPF406Obo+GEh1aOb/y3KYXz
9W5Qxdcv8wknG9UjD4TCE+icCz0OnRMY3uZ8iy/QNMgt6Wf8sQunwa0Ri4fjocO/kEkW+u4xaZ2s
pr44vbXlx3H+6XxlDlnis57kYFRbSwIBU/kc8Hs8DB4nDUogkfsrVZcNfqWzVrmdj0McpOmjIig5
+obeAtYDDtM0p/e0olNXk0RDfkmtsKViNbVfYRBrh9pEjC4/JL6djBwN9/r7q9F40iETlLbSVbnH
L54dK5Ef2wgosulp+x0DGf12r9qr6fQo7++rWOCaUQhLAMbqyFXz4NRGwz00xxNgnpn2cApZbitB
F2Vynmnep43EWWFi8fW3kXT+nAwoS1r/Xp1S/QxrLX2iNV57dVTkX1QZJi6eO1X4fP8IJP2ph7qr
MVziNdJQ3+ORCGkALVwkYMA8ArQeM9ErU4stgjyc+Uid/zXkXEbBW66v34ae5mKSY4+f/F1KmEbf
X/91o7t8lgJdx3so6wGd4tHYG9govLmZc4g8avR88Md2YmvUUJprZXfpuiodKCvbgVAtFpXO85Cz
DuCtvmloxWUcuJgIdOQY4uT8rB54THpMMEtOHVtZewLsBwvCTd+ONaBEAV4/X2HSViGhc0tAZklu
Cj1qcM4wWBu7UPvLQCi9G04xyoPU2hZm1MyaKCkynPZEqfcSLK20dZ5C2c74DkoxdMkuH6qxQhTh
ei7E3YQlULGU2aPPHa7hkrizM8ZerWExpVSDZI4rF/gQ1eHUI4mT9Uq55ZRMc5REjDox+Fb/HdZS
Pky5QYTbSKkikMiYEr3Uis6NGvy4tcdfhMfY8mcFpw+PbLqk+nkrb518zZ52Th6rbzspmPqqWUPU
Mf89Q2PFxXvs2/ngeEffrJHF0cTMCukDa6uFDcKUki29Xeax6EA+sxWYNaMa7nwFcxBPydpeQ7Fe
u3RJ6hoXViVWm+RxP0XcIlqLLJSlUqcDwkaQOWwoOfptvoFiLZ2b9nbBQI60XQgRPMG0zF4I5oKV
Rsi05LJenCUa1bHUcd3Yk4HLLpUVczhYt8xqsjlnI1VjycFknY0e+1Lhiu7iNh0stWbu8/QgHurA
JtIjCdR/ugrwpdfZWK5lmrGRgM83BF6D7ezU5StfadqPE/wvnt4w+zRgWH/altFGFnGBf9Qhqscj
eOy6HEmKlBkb7RV9q34wYb/mRGvGvvJ+eLs+SG3U5vLet8ASU0MO/ex4jq9wwZ7BOKHnQZtQk3Bb
DWN58CzarisCdyrFJ170663GdcFUav3QcO9FA2w8seapCLugYXsVSoL8eMexg/8Ge+eLkUANNAlR
CNnYdjzf9S3vA3wNCM7PwU7fFJa3WLyFFjGQRP+XVMBfKknmpUXMTiDUX4danYc8uNHzgyCVDFAd
EzhsSU7OzK7wEyDvTBv+v6vI60mKXFS8+/bsIFvUDenEjong/Tpb1LAnvI7xv7dnXRVMyLn0QhK3
ifvt2bd8M837KtwR6Er9qRQp9YWfYgQ0c5Lb/+q+v+sSg3hh6uUTspoDWbiDcJFdwWzyS/dLXpV5
CHQqf2CrvGGpm83eWy1690nQpiNiYqqfAsu8p+fGXBEMKCoPjctZ/BPD2xsq6H5IQrnL4/uR51hM
NQTTy7AP2iuOb98rgjUV9hBZ2J299e8+zWVVYND0CjYnDr/LqZweieixY2F9aCFf22+JSOhiV58H
MG+2Ixu5dN+jqxFj+iqAGEI//qWUgMDmxHuZqeYvn4Ag9/0osuM+CnIGHvsZmR7OOQLuGqr41ooG
akKEC56x4ZOxOLL3JUqh/MQpYeKicmn2II7+GHsdk3OYXmyR7kbc/ix/XJih9wsR6+fFfFNKc8VG
W8qtThvTmvr/aPr800BzoZ0/AbcWSN+TRsDjNaeT0u9hg66vZvUIUZgjGJSHI71f7mr72vCSPxnc
CC4eAiPGNQxFl3B+sJrv1SPvl24g/0bsVT+TbCuvjxOWmhCIFzg4Xg/gOAi61EmICy9irOA+iYUy
IE7761/Peo40yWuCU/IW4McDeIgV/namDpNa2WOLGShYkx27Di0hx+WHagK7Y4kswVlyBCub+BO6
JrbzWe2WRvNowLfxQTjh8RcSbcnboiwROO3aXdXYu3Q2h9iksK+UnvghmrExDo9yqb9Y9X1qcstU
a1GYFA0+oz06ZDENiEmUi0KZfO+LEXNmJ/srrYwOHuv+pfZggMH/rahO3YlQYscWiwSNqz4D3X82
+euamFvJ5vnRbFt/1TKGZ7hZGzTGesad0YOT/dls1q/8jK98BB5XgyJx8S+V4+TNT8m4N5D0dLdY
w79HQ1YYybQ9Ut1MtH/5Hmn+VK/FKSflje1zF/t2xC8nIgC+0rWQaReDaP2696DBdgxQWZEdCOgU
qYx/FAJm0kmaj3lWxopVNTlXaLx3HTqFf2wB6ah6vKbt3rXNANQpZAgaD7ELiC/aGGipryxeD98z
zIgOO5uZ3WzHCGObmDJQSbdaD2kSkPKcsPa7ATLFCuBHMjOSu1eQfMSjiMwe4V5gzriMJF0+erii
KJ5hh6XqZgKVPERW12tHTZFoOY+ISq+psGu2DWUTfiglfVfzFEuYrnZ/eaXgFFO8jOp/3g5Tcv8m
dtgE3kImwexjfpYcymLlSpi/uplUJFWrrIyFY0U2V3WToR6Lh+G70U4GtoPMO/iOwJl6png3In0r
cn/g1/4hdfVdVSEc9GnakWxM7gOtprM+Z/DsF/wacDvk9YezmzR3+mVzKlEhrZFNvvbbdv9sIiq2
RreOHn9rwDp8h/wWrSSmgxX88ZH65dVohihAun1rfC0RgJrSsxbFMhysZMsTB0Zs+5t9TwRq9GCz
WQDZ2d0DFwtdCmt2gJCgjKGTQNOpSuGxDnsmhA0/yX++JqFDuqXQQpw1023RfI17oyu4v6Yi16oY
KwVPymRv9kNJIjRg+CN6DNsBv3+4w856Z06eYN2zciT4xmpIf8uxNrnmZVW1qmtgAiN3+YgcfbUD
EebJbo4Pgt1shmZJ/zFdc+soWQ2hTlbEZR5dl4eyZgyeYKpKyXamFzWX3OhcpJ1hnFuxRAmWOr8/
NeP9RImcDlQDA0NP1EIzaXMfkDX4YVHEuguxMAcAKwErTZ+J/sQ220gWM21mNFnxhCkErLVl6/15
qPrDV+GzTWQITAXiRRumeStChuBoig14IeKcGiYLlX5qCr19tJ6RkCXYqTrM1jOhZ5cCWYDf1axb
oZA/cYNKdtVRZCmhPiO67YwA4y8KeYjxfWAaD56XnXzrbehpaI1ANnjuOB3wyrsB2EQNBzUn3i+8
TqzkFMLjPhb7vTyr8zlpnjf3NPkcZIXdN+YAep5/znE4oayX8aRJTKVLDcSm5ahVPPESpXvOyFBr
SsyP9tP6H82U/bDWQvmBKa/nNZHnhOrScIq9/Ia9/wukLp1PU9PTv+2EAvBasNrsDMROKOIgDdwO
tePHP2L7Lu2iH2yeDxbibUD1iLVb9kYKvFhLivXauSaSHlvcknAD+Prkiy8S6/CeYfK8pvcXijLn
MQdET/J+uyoePXOV7+kdm25QtkDEsq6YyfEu2zecN1uKclVqDtHb3ucPsuvOzobyo6X5Xk7HCDBd
1cb8N50ekdfTN+wga58JLS3vX2BN2p7PfMxofiAhDucb91kWePfT/GtPMb5/eDxMIAa8cugBKQYg
lr+DNFAzh97EJsKAOPzV7swnFOMUZco+4TgIU3utX9DNHw48jESZpvZSyVP7Y8Trssi3xaUUF+XU
g3ER2DjMXSmMXA/Rx4VDDdlBfc5/1FqjoVTYdITi1YtvpJ/DAKygcltYgiZu4/YXye+a79a5JPZ7
s2Ka4P3PBAJFo/GOFW1Jy6dkRltpFAn/txY1QPPKoGZsEy9fgSU5e3QO+cbKyfRWZs1Glg3NLNK7
1qWIS3B+EqtJiI7Ges+h5rKvjVHtoH+RSoVVaBker3N/vXaJGgcIk+pRiPmqiBlX+ypJD/MRgt5h
TnixZiUp8eOQKITNtvI83n0Qmf2dGGeLkZyqsome7jY4ZekP+/BrKblsB922YmSBAPzHyfEZzVzr
/Xydy49WUY09eh9isZtObfQ/Sg1Tz/udtEeM/YbYb/sMyoaFjxorbwVLd9FRD725uWU65o6LnrIG
xrXFUnTdfRXbk13j6oxsqRwC+TdWWnK+fFUhvZnErcNLUT/ZXHq+kptRY7D52p+iXPjXYOf8v5Bk
kbyKrHP1x9Qib7a9R3qbBxiZucwlCAPCzHjUYojAZUeyC3Vt6wY21dzmqCChqoBEP49hn47N64Yw
y6lKYsBzIRBnPvVZcvmhWBDSVngagvlIrBR/0mFlx3NQn0+SQ8Jh6ZYMR/DozkbBIkOSdOAIYN2x
jhTM4TMFLEtwCE/WT+v0gC9z00c0/upNq8lBroTg9dJsN83RGjKiwzCnEbjxPrrJ9pgh72u4ZC6f
nbCrtHE5gI7EdYFI0HdHlPv3QrA2p7+eRB/z1MM+qpg7FZmLhMRO4GYAd3eqAqkyNV09Zf9yb4EZ
mYF9pj0dBOJtKlR2Zj4QrHUOnalZ0kS4mJl03bZ2jjnhRRUezGHfcECSsaUq5CKJIPuiUm3eCJBo
BeVf2UQhzPCNsSNZWhkmVo9h5bYamqmiyrKZHcPF7LFS/65XHAPfR1IMwRQqnL2csM7971cZDCkY
fd8a5L6Z6mi1RysyJ7kdHqweNUq9/YVBdBqYVzKXnjfyE15t3BPd2+0rXrQqQmOV+RrBEJ88vXPO
uRoDpLHYzyoHKhKew4u+9aA1h75klM/NXiHbV7i0CQhyLA5ClSGc7ht6YIQNYpeUfP6z/WqOVOB8
LYN8NuKW7rY5vAUpi/vzEus/1kGDskJLyCuF6mEDUO1iBYF7Fs+56fwm0Y5OgEfq6Gerq5x8iw7n
v4EW+y1wqjBc+EjxPGU9OJvYaFi7jkpu1MR3vmuwQLTzyhXjl3I2pXnc9QteGrLfr3jKpmYMOzcj
j7hFfvcQ3HhkY7xmvVTYYxg6KWWeFtkyiK6QkyIM0Lqdwe6DOs3dVEO0ePNnk6dYyt3biDLX3HMr
YJdLXj2M7/bEBgOE2d+GLnAggi7bWlO2onTndd38KNlzTm7n1SACSEMwZ9WMAKaA1iVewTZmb/aY
MofNpTl0qO9ks+0QBwk6P8VFQKpTu+roP1S5rNpHBZ6SIq/yyrwpoe7Q5h3dbFGWl2sIJHIdKUjm
rIiGyRBL96BbZo09vGkn88NVyWgdiVeszkeweDx3P9mSEf1lNlY+w5sgmTbQX2oS+tlTRRKzFnyU
1K4PYlSekk9aIPrzBzLlm6Oi606WPJBHEhPvzvsJZAW/74/CcmT75XoXrM8SvUpK4ZSS0I7xkl25
lpEiez/39HsJjq9jzrLpY6K/oPHZdbEhHBwf5X/GJX4BUyChQ1UNyoa0dJi1t209N+vu9Wt3noqC
pnsCnz//mrLBYkIyGmTZrTqubAf/FZqu+emNPHz3hX/592KLF1cB33d9addTl5O/I2TSSd+wkRli
Y+mUKKtzWHvQe5VUgfSPSQVxWH6yYC+HTxb+6E5M1wMmT0QBzuHDekZQ9hugjsxfPq9veaLB7syy
GPoAfiigy+Qi6ra+uYTK1+XnzkqEhMKb6oBdFzmVGlEGJtjuxWOuwDjXgAtFoBSuCDBaQcmZNGws
n8HjlG72G/g9HJzHdk1YyUjGSnU1xL9tw43Fn2RAA00jSJTWjlKiviS0v+nSWo8uiJX+wNFG8XZe
kUHlwLKLBL0/Vvg/QIcOvWgnbTRL8z6RnYrC1eqz+ObG9yhQKllOslNCLDbxvkoeXK2/YtLj5EdR
GpVfRxGfdPYgpJXgRFwdFhBfWXlAsjUEsh8elNsxaUNuvadTbD+HsWUnNHyVHk6dQnzhBOY4DwBE
nOkXvEiHz1nF/rCUuTrr7ch6+DxHMyHN4frGQv7quSUprmbdY6mgiLdFlOnvGf3d5co0dY/306d3
3YluD9qrZJosocw6/LektsJUz0gUvixwECnEsxKCfW4T13KtrAJ/ODSIKEkB4hJT5DPVTQa63GbD
lCM6QuXMPC+SpPVq03AUyBu497Xyi6iiyy7sPmOSeCSBmRyPSX95PBpsqgeNdUJXJ9+KQKe7jhev
kKCsmMI1OUrwp2U8mExGJ54HB6N7cYI2x+XW0K5Lq3/SOsbtsidJcH6GYPF4nbvdE+X7y8A2I7hd
FVLby/2+7NNhdA+b7F5FS+aD8JNaHZ/Hb253nYfFrowXulgkD+XX/yE2skYA2emECktN3bKGaFOi
zOrL4JwwRX71yTP0eTYtefkGkimG17UTeQCZjECLKSWoKPqQlR3Fg64E5SRN+tPKv4Zjp1CYqq4e
Y7BpMcLojc1g7pER4ENm0uxGer0eiObQ9yvqNvmwLBDHD3cbBkYZEOYVxHh/vyyyesMK9VYKPQiH
YzVIWb4tc189DKWWpUVmCVNLUN5wLaC90gbfvDfyGwG1wbaHQqYtXf3p7FJ/rNhXtXGg+3NceJXd
+HxkNU7T+0bBqVAylXfgavYGXInCXdx/8Z8lsIZiOe9kSLiaS5asGCRp8QGvjyroQ2bShb4SEYxX
BfOQbGnUcNxmmxbkfr2z8z8JQZPfFYpJQIuSv42BvmWJPKJOquLyeh4c50lwmhjHUX0XC3SoUEBw
z5AwVOBcAhQEBtE/ufxS+P4nZM/+rqStkw7UG0/eoKs2IeDQMzXE/0vZ4rpgVCkbYH1hggFeKNZ8
5bzCwXGNem6HeCKs77Y0p/+5Rf1v+de1wcKnYb+g+Zyz6GX724+YIpnb302w5huRhvI99SzZY0pB
8Q==
`pragma protect end_protected
